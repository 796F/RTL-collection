-- =====================================================================
-- Copyright � 2010 by Cryptographic Engineering Research Group (CERG),
-- ECE Department, George Mason University
-- Fairfax, VA, U.S.A.
-- =====================================================================

library ieee;
use ieee.std_logic_1164.all;

package sha3_hamsi_512cons is
	type gen512_type is array (0 to 31, 0 to 255) of integer range 0 to 3;
	constant generator512 : gen512_type := (
		(1,0,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,1,2,2,0,1,2,3,3,2,0,0,2,1,3,3,2,1,1,0,2,0,2,1,1,3,2,2,1,3,0,3,2,3,2,0,1,1,0,2,2,0,3,0,0,3,2,2,2,0,1,1,2,0,0,2,1,2,1,0,2,0,3,0,
		3,2,3,1,3,2,1,2,2,1,2,0,1,0,1,0,3,3,1,0,1,0,0,1,3,3,1,3,3,1,2,2,3,1,3,2,1,2,3,3,2,0,0,2,1,3,0,3,0,1,3,1,3,2,1,2,1,2,2,1,0,0,1,0,0,1,3,
		3,1,3,2,2,1,3,3,3,1,2,2,1,2,2,2,2,2,2,3,1,3,2,1,2,1,3,3,1,2,2,3,3,3,3,3,3,0,3,0,2,3,2,3,2,1,1,3,2,1,3,0,3,0,1),
		(0,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,1,1,0,2,2,0,0,1,3,3,1,2,0,2,3,0,3,2,0,0,2,1,1,1,0,1,2,0,2,2,1,2,0,1,0,2,1,1,2,3,3,2,3,2,1,3,1,2,1,3,3,2,1,1,3,1,0,3,0,3,0,0,3,
		2,2,1,1,1,1,1,1,1,3,0,3,0,1,1,3,2,2,1,3,3,1,3,2,1,2,2,3,3,2,0,0,1,1,1,1,1,1,0,2,0,1,2,1,0,1,2,2,0,1,1,1,1,1,1,1,0,0,3,2,2,3,3,1,3,2,1,
		2,1,0,1,2,0,2,2,0,1,1,2,0,2,3,1,3,1,2,1,1,1,1,1,1,2,3,3,2,0,0,3,1,2,1,2,3,3,0,1,0,1,3,3,0,3,1,0,1,0,1,2,2,0,1),
		(0,0,0,0,1,0,0,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,2,3,2,1,3,1,1,3,3,1,2,2,1,0,1,2,0,2,0,2,3,3,0,2,2,1,0,1,0,2,3,2,1,1,3,2,0,1,2,2,0,1,3,3,2,0,0,2,3,3,0,1,1,0,1,1,1,1,1,1,3,3,2,0,
		0,2,2,2,0,3,3,0,1,1,3,0,0,3,0,2,0,1,2,1,2,0,1,1,2,0,3,2,2,3,1,1,3,1,2,1,2,3,1,0,0,1,3,3,1,3,0,3,0,1,3,3,1,2,2,1,3,0,0,3,2,2,1,0,1,2,0,
		2,2,3,3,2,0,0,0,2,3,3,0,2,2,1,0,1,0,2,0,1,2,2,0,1,1,0,2,0,2,1,0,2,0,1,2,1,3,0,1,0,1,3,1,2,3,2,3,1,3,1,1,3,0,0),
		(0,0,0,0,0,1,0,3,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,3,0,1,0,1,3,1,2,0,0,1,2,2,0,1,1,2,0,1,3,1,0,3,0,0,2,1,2,1,0,2,2,3,1,1,3,3,2,3,0,2,0,3,1,1,3,0,0,0,3,3,0,1,1,2,0,0,2,1,1,3,1,1,3,
		0,0,0,2,2,0,3,3,1,2,2,1,0,0,0,0,2,1,1,2,2,3,1,3,1,2,3,1,0,0,3,1,3,1,3,2,1,2,0,1,0,3,1,3,0,1,3,1,3,0,2,2,2,2,2,2,0,3,0,2,3,2,2,0,1,1,2,
		0,1,1,0,2,2,0,1,3,1,0,3,0,0,2,1,2,1,0,3,2,3,0,2,0,3,3,2,0,0,2,0,0,2,1,1,2,2,2,1,0,0,1,1,2,1,3,2,3,2,2,0,3,3,0),
		(0,0,0,0,0,0,1,3,3,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,2,2,1,0,0,1,0,1,2,2,0,1,2,3,1,3,1,2,2,0,2,3,0,3,2,1,3,3,2,1,1,1,1,1,1,1,1,0,1,2,0,2,2,2,0,3,3,0,1,3,0,3,0,1,0,2,0,1,2,1,2,2,0,3,
		3,0,3,2,0,2,0,3,3,3,0,1,1,0,3,2,2,3,1,1,2,3,2,1,3,1,0,3,1,1,0,3,1,0,2,0,2,1,0,0,1,3,3,1,1,3,2,2,1,3,3,0,0,3,2,2,0,0,3,2,2,3,2,3,1,3,1,
		2,0,1,1,0,2,2,2,0,2,3,0,3,2,1,3,3,2,1,1,0,1,2,0,2,3,1,1,3,0,0,3,2,2,3,1,1,2,3,3,2,0,0,2,0,3,0,3,2,0,2,2,0,3,3),
		(0,0,0,0,0,0,0,0,0,0,1,0,0,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,2,2,1,0,0,1,2,0,1,1,2,0,1,3,2,2,1,3,0,1,1,0,2,2,2,3,2,1,3,1,1,3,0,3,0,1,3,2,3,0,2,0,2,1,1,2,3,3,0,2,3,3,0,2,0,2,3,3,0,2,0,3,3,0,
		1,1,0,1,1,0,2,2,1,3,0,3,0,1,3,0,3,1,0,1,0,3,0,2,3,2,1,0,2,0,2,1,2,3,1,3,1,2,3,3,3,3,3,3,3,1,0,0,3,1,3,3,1,2,2,1,3,1,2,1,2,3,0,1,1,0,2,
		2,2,2,2,2,2,2,2,0,0,2,1,1,0,0,2,1,1,2,0,1,0,3,1,3,3,2,3,0,2,0,2,3,1,3,1,2,3,1,1,3,0,0,3,3,1,2,2,1,2,3,2,1,3,1),
		(0,0,0,0,0,0,0,0,0,0,0,1,0,3,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,2,3,3,2,0,0,2,3,1,3,1,2,3,3,1,2,2,1,2,1,0,1,0,2,3,0,1,0,1,3,0,1,3,1,3,0,1,0,1,2,0,2,2,3,0,0,2,3,1,3,1,0,3,0,1,3,1,0,3,0,1,3,0,3,
		0,1,2,1,0,1,0,2,0,1,3,1,3,0,1,0,3,3,1,0,0,0,3,2,2,3,3,3,2,0,0,2,2,3,2,1,3,1,1,0,0,1,3,3,0,3,1,1,0,3,2,2,2,2,2,2,3,1,3,2,1,2,2,1,0,1,0,
		2,3,0,0,3,2,2,0,2,0,1,2,1,3,2,2,3,1,1,0,0,1,3,3,1,1,0,1,2,0,2,2,3,2,1,3,1,2,2,0,3,3,0,2,2,2,2,2,2,3,0,1,0,1,3),
		(0,0,0,0,0,0,0,0,0,0,0,0,1,3,3,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,1,1,0,2,2,0,2,3,2,1,3,1,2,2,2,2,2,2,0,2,1,2,1,0,2,2,1,0,0,1,1,3,2,2,1,3,2,0,1,1,2,0,0,2,3,3,0,2,2,0,2,3,0,3,2,0,2,3,0,3,0,1,3,1,
		3,0,0,2,1,2,1,0,1,3,2,2,1,3,1,2,3,2,3,1,1,3,3,1,2,2,3,1,1,3,0,0,3,0,1,0,1,3,0,1,0,3,1,3,2,1,2,0,1,0,3,0,0,3,2,2,1,0,2,0,2,1,0,2,1,2,1,
		0,0,3,0,2,3,2,0,0,2,1,1,2,3,1,0,0,3,1,2,1,1,2,3,3,2,0,1,1,2,0,3,0,1,0,1,3,0,2,2,0,3,3,3,0,0,3,2,2,2,2,1,0,0,1),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,1,0,3,1,3,3,0,1,0,1,3,1,3,3,1,2,2,3,2,3,0,2,0,3,0,0,3,2,2,2,0,3,0,3,2,0,2,3,3,0,2,0,2,3,3,0,2,2,1,3,3,2,1,1,3,2,2,1,3,0,2,0,1,
		2,1,2,2,3,1,1,3,3,2,1,1,3,2,1,1,3,0,0,3,2,0,1,1,2,0,0,2,3,3,0,2,1,3,2,2,1,3,3,0,0,3,2,2,3,1,0,0,3,1,1,0,3,3,1,0,3,1,3,2,1,2,3,1,0,0,3,
		1,2,0,1,1,2,0,3,0,2,2,3,0,3,3,1,2,2,1,1,2,3,2,3,1,2,1,1,2,3,3,0,3,1,1,0,3,0,3,0,2,3,2,0,1,0,3,1,3,1,0,3,3,1,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,3,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,1,3,3,1,2,2,1,0,0,1,1,2,0,0,1,2,1,0,1,2,0,2,0,3,0,2,3,2,1,1,3,0,0,3,1,3,1,0,3,0,1,3,1,0,3,0,1,1,2,3,3,2,3,3,1,2,2,1,0,0,2,1,
		1,2,1,1,1,1,1,1,2,2,3,1,1,3,1,2,2,1,0,0,2,3,1,3,1,2,1,3,1,0,3,0,3,3,1,2,2,1,0,3,0,2,3,2,0,3,1,1,0,3,1,2,3,2,3,1,1,0,2,0,2,1,0,3,1,1,0,
		3,2,3,1,3,1,2,3,1,2,1,2,3,2,2,2,2,2,2,1,2,1,3,2,3,2,3,0,0,2,3,2,1,2,0,1,0,0,0,3,2,2,3,0,0,1,3,3,1,1,2,3,2,3,1),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,3,3,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,2,1,1,2,3,3,2,3,3,2,0,0,0,1,2,2,0,1,2,0,1,1,2,0,0,0,3,2,2,3,1,2,2,1,0,0,2,0,2,3,0,3,2,0,2,3,0,3,3,3,3,3,3,3,2,2,2,2,2,2,3,2,2,3,
		1,1,2,0,0,2,1,1,1,1,1,1,1,1,3,3,0,1,1,0,2,3,2,1,3,1,2,0,2,3,0,3,2,2,2,2,2,2,0,0,3,2,2,3,2,1,2,0,1,0,1,2,1,3,2,3,3,3,2,0,0,2,2,1,2,0,1,
		0,2,3,2,1,3,1,3,1,3,2,1,2,3,0,0,3,2,2,2,0,3,0,3,2,0,2,3,3,0,2,3,0,3,1,0,1,1,3,3,1,2,2,2,1,1,2,3,3,1,2,1,3,2,3),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,3,1,0,0,3,1,2,1,2,0,1,0,3,3,2,0,0,2,3,2,1,1,3,2,2,1,3,3,2,1,1,0,1,2,0,2,2,1,2,0,1,0,2,3,2,1,3,1,0,3,1,1,0,3,2,1,0,1,0,2,1,1,1,1,
		1,1,2,0,3,0,3,2,2,0,2,3,0,3,2,2,2,2,2,2,2,2,3,1,1,3,1,3,2,2,1,3,2,1,3,3,2,1,0,1,1,0,2,2,2,0,3,0,3,2,1,1,0,2,2,0,0,3,1,1,0,3,3,0,1,0,1,
		3,1,3,3,1,2,2,0,0,3,2,2,3,2,2,1,0,0,1,1,0,2,0,2,1,0,2,1,2,1,0,3,0,2,2,3,0,1,3,3,1,2,2,2,1,0,1,0,2,1,1,3,0,0,3),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,3,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,3,1,1,0,3,3,0,3,1,0,1,3,1,1,3,0,0,2,2,3,1,1,3,1,1,2,3,3,2,2,0,1,1,2,0,3,0,3,1,0,1,3,0,1,0,1,3,2,1,2,0,1,0,0,2,1,2,1,0,2,0,0,2,
		1,1,1,1,3,0,0,3,3,0,2,2,3,0,3,0,0,3,2,2,1,1,1,1,1,1,3,3,1,2,2,1,1,1,2,3,3,2,2,1,0,1,0,2,1,1,3,0,0,3,0,1,1,0,2,2,2,1,2,0,1,0,2,2,1,0,0,
		1,1,2,0,0,1,2,1,3,3,1,2,2,2,3,3,2,0,0,3,3,2,0,0,2,2,1,3,3,2,1,3,1,2,1,2,3,1,2,0,0,1,2,0,2,1,2,1,0,1,2,2,1,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,3,3,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,2,1,2,0,1,0,1,0,3,3,1,0,2,2,0,3,3,0,1,1,1,1,1,1,3,3,3,3,3,3,2,3,1,3,1,2,1,0,3,3,1,0,2,2,1,0,0,1,3,0,3,1,0,1,2,1,3,3,2,1,0,2,0,1,
		2,1,1,2,2,1,0,0,3,1,2,1,2,3,0,3,0,2,3,2,2,0,0,2,1,1,2,2,2,2,2,2,3,3,3,3,3,3,0,2,1,2,1,0,1,2,2,1,0,0,2,1,0,1,0,2,3,0,3,1,0,1,2,3,3,2,0,
		0,0,1,2,2,0,1,1,2,0,0,1,2,1,1,0,2,2,0,3,1,1,3,0,0,1,1,2,3,3,2,3,1,3,2,1,2,0,1,2,2,0,1,2,1,3,3,2,1,3,3,0,1,1,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,2,2,3,1,1,3,3,0,0,3,2,2,3,3,1,2,2,1,1,3,2,2,1,3,2,0,0,2,1,1,2,1,0,1,0,2,3,3,0,1,1,0,0,0,1,3,3,1,0,1,0,3,1,3,0,2,2,0,3,3,1,2,3,2,
		3,1,2,0,0,2,1,1,1,0,2,0,2,1,2,0,0,2,1,1,3,2,1,1,3,2,3,3,3,3,3,3,0,2,0,1,2,1,1,3,1,0,3,0,0,1,3,1,3,0,2,2,1,0,0,1,0,0,3,2,2,3,2,1,3,3,2,
		1,0,1,0,3,1,3,1,2,3,2,3,1,3,2,1,1,3,2,3,2,0,2,0,3,1,2,1,3,2,3,2,3,3,2,0,0,3,2,1,1,3,2,2,3,1,3,1,2,3,0,3,1,0,1),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,3,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,1,1,1,1,1,1,0,3,0,2,3,2,2,2,2,2,2,2,3,3,1,2,2,1,0,2,0,1,2,1,0,2,1,2,1,0,0,3,3,0,1,1,2,1,1,2,3,3,0,0,1,3,3,1,3,2,0,2,0,3,1,2,1,3,
		2,3,0,2,0,1,2,1,3,3,2,0,0,2,0,2,0,1,2,1,2,2,3,1,1,3,1,0,0,1,3,3,0,0,2,1,1,2,2,0,2,3,0,3,1,3,2,2,1,3,2,3,3,2,0,0,1,3,3,1,2,2,1,1,2,3,3,
		2,0,0,1,3,3,1,1,2,1,3,2,3,2,2,3,1,1,3,0,3,2,3,2,0,2,0,3,0,3,2,1,1,0,2,2,0,2,2,3,1,1,3,2,3,2,1,3,1,1,0,3,3,1,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,3,3,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,2,0,0,2,1,1,0,0,3,2,2,3,3,0,0,3,2,2,2,2,2,2,2,2,0,0,2,1,1,2,2,1,3,3,2,1,1,3,0,3,0,1,2,3,0,0,2,3,2,1,1,2,3,3,0,3,2,3,2,0,2,0,3,0,
		3,2,0,0,2,1,1,2,3,1,1,3,0,0,0,0,2,1,1,2,1,1,1,1,1,1,0,1,0,3,1,3,3,2,2,3,1,1,3,0,2,2,3,0,3,3,1,2,2,1,1,1,0,2,2,0,1,2,0,0,1,2,3,3,3,3,3,
		3,2,1,1,2,3,3,2,0,3,0,3,2,1,1,1,1,1,1,3,2,1,1,3,2,1,1,3,0,0,3,0,1,1,0,2,2,1,1,1,1,1,1,3,0,1,0,1,3,1,2,3,2,3,1),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,3,3,2,0,0,2,2,3,2,1,3,1,3,0,2,2,3,0,1,1,1,1,1,1,2,1,0,1,0,2,3,3,0,1,1,0,2,1,3,3,2,1,0,3,1,1,0,3,1,2,3,2,3,1,1,3,1,0,3,0,2,1,1,2,
		3,3,0,1,2,2,0,1,3,2,0,2,0,3,2,2,2,2,2,2,2,2,0,3,3,0,2,2,0,3,3,0,1,1,2,3,3,2,0,1,2,2,0,1,2,1,1,2,3,3,3,1,1,3,0,0,2,1,0,1,0,2,1,2,1,3,2,
		3,3,2,2,3,1,1,0,0,1,3,3,1,1,1,1,1,1,1,0,2,1,2,1,0,2,3,2,1,3,1,0,3,0,2,3,2,3,2,1,1,3,2,3,3,1,2,2,1,1,3,2,2,1,3),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,3,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,3,1,1,3,0,0,3,0,1,0,1,3,3,1,2,1,2,3,2,0,0,2,1,1,0,2,1,2,1,0,0,3,3,0,1,1,1,1,2,3,3,2,2,1,2,0,1,0,1,2,1,3,2,3,2,0,2,3,0,3,2,3,0,0,
		2,3,3,2,3,0,2,0,0,3,2,3,2,0,3,0,0,3,2,2,0,2,2,0,3,3,0,2,2,0,3,3,3,3,3,3,3,3,3,2,3,0,2,0,2,3,0,0,2,3,2,2,0,3,3,0,0,2,1,2,1,0,2,0,3,0,3,
		2,3,1,0,0,3,1,2,1,1,2,3,3,2,0,0,2,1,1,2,1,3,3,2,1,3,0,1,0,1,3,0,0,3,2,2,3,2,2,3,1,1,3,2,2,2,2,2,2,3,3,1,2,2,1),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,3,3,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,2,2,0,3,3,0,2,2,1,0,0,1,3,1,3,2,1,2,0,2,0,1,2,1,2,1,3,3,2,1,1,3,0,3,0,1,3,3,3,3,3,3,3,0,3,1,0,1,2,0,3,0,3,2,3,0,2,2,3,0,0,2,3,3,
		0,2,1,0,1,2,0,2,3,2,1,1,3,2,0,3,0,2,3,2,3,2,0,2,0,3,3,2,0,2,0,3,1,0,0,1,3,3,1,0,1,2,0,2,0,2,3,3,0,2,0,2,2,0,3,3,2,1,3,3,2,1,1,1,3,0,0,
		3,0,3,1,1,0,3,2,3,0,0,2,3,0,2,0,1,2,1,1,1,2,3,3,2,2,2,1,0,0,1,1,3,3,1,2,2,1,1,1,1,1,1,3,0,0,3,2,2,2,2,2,2,2,2),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,1,0,3,1,3,2,1,2,0,1,0,1,0,0,1,3,3,1,1,3,0,0,3,2,0,0,2,1,1,2,2,1,0,0,1,2,2,3,1,1,3,1,1,3,0,0,3,0,3,3,0,1,1,0,3,2,3,2,0,1,3,2,2,
		1,3,0,0,1,3,3,1,3,2,2,3,1,1,3,0,3,1,0,1,3,2,0,2,0,3,2,3,3,2,0,0,2,1,0,1,0,2,0,2,3,3,0,2,0,3,1,1,0,3,0,0,2,1,1,2,3,3,3,3,3,3,2,1,2,0,1,
		0,3,3,1,2,2,1,2,0,2,3,0,3,1,3,0,3,0,1,0,3,0,2,3,2,2,2,0,3,3,0,1,2,0,0,1,2,2,3,1,3,1,2,0,2,0,1,2,1,2,0,3,0,3,2),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,3,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,0,1,3,3,1,3,0,3,1,0,1,0,1,0,3,1,3,1,2,2,1,0,0,0,2,0,1,2,1,2,3,3,2,0,0,1,1,1,1,1,1,1,2,2,1,0,0,1,3,0,3,0,1,3,2,1,1,3,2,3,3,1,2,
		2,1,2,1,1,2,3,3,3,1,0,0,3,1,1,0,3,3,1,0,0,3,2,3,2,0,1,1,0,2,2,0,0,2,1,2,1,0,1,3,1,0,3,0,2,1,2,0,1,0,3,2,2,3,1,1,1,0,0,1,3,3,3,0,3,1,0,
		1,2,2,2,2,2,2,3,0,2,2,3,0,0,1,3,1,3,0,0,0,3,2,2,3,0,2,2,0,3,3,0,1,2,2,0,1,2,3,2,1,3,1,0,0,2,1,1,2,1,1,3,0,0,3),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,3,3,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,2,1,1,2,3,3,1,0,3,3,1,0,0,0,1,3,3,1,3,3,0,1,1,0,0,0,2,1,1,2,1,1,0,2,2,0,2,0,0,2,1,1,3,3,0,1,1,0,0,1,3,1,3,0,2,2,3,1,1,3,2,2,2,2,
		2,2,2,3,0,0,2,3,0,3,1,1,0,3,1,2,3,2,3,1,3,2,1,1,3,2,0,1,1,0,2,2,2,1,3,3,2,1,2,0,2,3,0,3,3,0,3,1,0,1,3,1,0,0,3,1,0,1,0,3,1,3,1,0,3,3,1,
		0,3,0,0,3,2,2,3,1,2,1,2,3,1,3,2,2,1,3,1,3,3,1,2,2,3,2,0,2,0,3,3,2,3,0,2,0,3,0,1,0,1,3,3,2,2,3,1,1,1,2,2,1,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,1,2,0,0,1,2,3,1,3,2,1,2,2,0,3,0,3,2,2,2,3,1,1,3,3,0,3,1,0,1,1,0,2,0,2,1,2,0,3,0,3,2,1,0,1,2,0,2,1,3,0,3,0,1,0,3,2,3,2,0,0,0,3,2,
		2,3,2,0,3,0,3,2,0,3,3,0,1,1,1,2,3,2,3,1,2,1,3,3,2,1,2,3,1,3,1,2,1,2,3,2,3,1,0,2,1,2,1,0,2,2,2,2,2,2,3,3,1,2,2,1,2,1,1,2,3,3,3,1,0,0,3,
		1,1,2,3,2,3,1,0,3,2,3,2,0,0,3,3,0,1,1,2,2,1,0,0,1,2,3,3,2,0,0,0,0,1,3,3,1,3,2,3,0,2,0,1,0,1,2,0,2,2,2,3,1,1,3),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,3,1,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,0,1,2,2,0,1,1,0,2,0,2,1,1,1,3,0,0,3,1,1,1,1,1,1,1,0,3,3,1,0,3,3,2,0,0,2,1,1,3,0,0,3,2,0,1,1,2,0,0,1,3,1,3,0,3,2,1,1,3,2,1,3,3,1,
		2,2,1,1,3,0,0,3,1,3,0,3,0,1,1,2,1,3,2,3,1,1,2,3,3,2,2,3,2,1,3,1,1,2,1,3,2,3,2,1,3,3,2,1,3,0,0,3,2,2,2,2,2,2,2,2,2,3,0,0,2,3,0,3,1,1,0,
		3,1,2,1,3,2,3,3,2,1,1,3,2,1,3,0,3,0,1,2,3,3,2,0,0,1,1,0,2,2,0,2,1,1,2,3,3,1,0,1,2,0,2,2,0,1,1,2,0,1,1,1,1,1,1),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,3,3,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
		0,0,0,3,2,3,0,2,0,3,3,2,0,0,2,1,2,2,1,0,0,2,0,0,2,1,1,1,2,3,2,3,1,3,1,1,3,0,0,1,2,2,1,0,0,2,3,1,3,1,2,1,3,2,2,1,3,2,2,3,1,1,3,1,2,0,0,
		1,2,1,2,2,1,0,0,0,1,3,1,3,0,2,0,3,0,3,2,3,3,3,3,3,3,3,0,1,0,1,3,2,0,3,0,3,2,1,1,2,3,3,2,0,3,0,2,3,2,3,0,0,3,2,2,0,2,3,3,0,2,2,1,2,0,1,
		0,2,0,3,0,3,2,2,2,3,1,1,3,0,1,3,1,3,0,1,1,0,2,2,0,0,1,1,0,2,2,2,3,0,0,2,3,2,0,1,1,2,0,2,3,1,3,1,2,2,0,0,2,1,1),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,3,3,0,0,0,0,0,0,0,0,0,
		0,0,0,3,1,3,2,1,2,3,1,3,2,1,2,1,1,3,0,0,3,1,3,1,0,3,0,2,0,3,0,3,2,0,3,3,0,1,1,2,0,2,3,0,3,0,3,2,3,2,0,3,0,2,2,3,0,0,3,3,0,1,1,3,3,3,3,
		3,3,2,3,3,2,0,0,2,0,0,2,1,1,2,1,3,3,2,1,0,3,2,3,2,0,2,0,1,1,2,0,0,0,3,2,2,3,1,0,1,2,0,2,2,0,1,1,2,0,3,1,3,2,1,2,0,1,3,1,3,0,0,1,2,2,0,
		1,1,2,0,0,1,2,3,1,0,0,3,1,0,1,0,3,1,3,3,0,2,2,3,0,2,0,0,2,1,1,1,1,2,3,3,2,0,2,0,1,2,1,0,1,0,3,1,3,3,2,2,3,1,1),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,3,1,3,0,0,0,0,0,0,0,0,0,
		0,0,0,1,0,2,0,2,1,1,0,2,0,2,1,1,2,2,1,0,0,2,0,2,3,0,3,1,1,3,0,0,3,1,3,0,3,0,1,3,0,2,2,3,0,3,2,1,1,3,2,3,1,2,1,2,3,1,3,0,3,0,1,1,0,0,1,
		3,3,1,1,0,2,2,0,0,2,0,1,2,1,1,1,2,3,3,2,3,2,1,1,3,2,2,3,1,3,1,2,1,3,3,1,2,2,2,0,1,1,2,0,2,3,1,3,1,2,1,0,2,0,2,1,1,3,2,2,1,3,3,2,3,0,2,
		0,0,1,2,2,0,1,0,3,1,1,0,3,0,0,1,3,3,1,3,1,2,1,2,3,0,2,0,1,2,1,3,3,3,3,3,3,0,0,2,1,1,2,0,0,1,3,3,1,3,1,0,0,3,1),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,3,3,1,0,0,0,0,0,0,0,0,0,
		0,0,0,3,3,2,0,0,2,3,3,2,0,0,2,3,3,0,1,1,0,3,0,2,2,3,0,1,2,2,1,0,0,0,1,3,1,3,0,3,1,2,1,2,3,2,2,3,1,1,3,3,1,3,2,1,2,0,1,3,1,3,0,0,1,0,3,
		1,3,0,1,1,0,2,2,0,0,2,1,1,2,3,3,3,3,3,3,2,2,3,1,1,3,2,3,2,1,3,1,1,2,0,0,1,2,2,3,1,3,1,2,2,3,2,1,3,1,3,3,2,0,0,2,3,3,1,2,2,1,1,0,1,2,0,
		2,3,2,3,0,2,0,2,1,2,0,1,0,2,1,1,2,3,3,3,1,3,2,1,2,0,0,2,1,1,2,1,0,0,1,3,3,3,2,2,3,1,1,2,1,1,2,3,3,0,3,1,1,0,3),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,3,3,0,0,0,
		0,0,0,3,1,0,0,3,1,1,1,1,1,1,1,3,2,0,2,0,3,3,0,1,0,1,3,0,0,1,3,3,1,0,0,2,1,1,2,0,2,2,0,3,3,0,1,3,1,3,0,0,2,0,1,2,1,3,0,1,0,1,3,0,1,0,3,
		1,3,1,1,0,2,2,0,2,1,2,0,1,0,3,0,3,1,0,1,1,2,3,2,3,1,3,0,1,0,1,3,0,3,1,1,0,3,1,2,0,0,1,2,0,0,2,1,1,2,0,0,1,3,3,1,2,2,1,0,0,1,0,0,1,3,3,
		1,2,3,1,3,1,2,3,2,2,3,1,1,2,3,3,2,0,0,2,2,3,1,1,3,2,0,0,2,1,1,3,1,3,2,1,2,0,1,0,3,1,3,2,0,0,2,1,1,3,3,2,0,0,2),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,3,1,3,0,0,0,
		0,0,0,0,3,1,1,0,3,2,0,0,2,1,1,0,3,2,3,2,0,2,2,1,0,0,1,2,1,1,2,3,3,3,2,2,3,1,1,3,2,0,2,0,3,1,3,2,2,1,3,0,0,2,1,1,2,2,2,1,0,0,1,0,0,1,3,
		3,1,0,1,1,0,2,2,3,0,3,1,0,1,1,0,3,3,1,0,1,2,1,3,2,3,2,2,1,0,0,1,2,1,2,0,1,0,0,1,2,2,0,1,3,2,2,3,1,1,2,1,1,2,3,3,2,3,3,2,0,0,2,1,1,2,3,
		3,2,3,2,1,3,1,3,1,0,0,3,1,1,1,0,2,2,0,1,1,1,1,1,1,0,2,0,1,2,1,1,0,2,0,2,1,0,0,1,3,3,1,0,2,0,1,2,1,3,1,1,3,0,0),
		(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,3,3,1,0,0,0,
		0,0,0,2,1,2,0,1,0,0,2,0,1,2,1,3,2,1,1,3,2,2,3,3,2,0,0,2,3,0,0,2,3,3,1,0,0,3,1,0,3,2,3,2,0,3,3,1,2,2,1,3,2,2,3,1,1,2,3,3,2,0,0,2,1,1,2,
		3,3,2,1,0,1,0,2,1,0,3,3,1,0,1,2,3,2,3,1,2,0,3,0,3,2,2,3,3,2,0,0,3,0,3,1,0,1,3,2,3,0,2,0,3,1,0,0,3,1,2,3,0,0,2,3,1,1,0,2,2,0,2,3,0,0,2,
		3,3,0,1,0,1,3,0,3,1,1,0,3,0,1,1,0,2,2,2,0,0,2,1,1,0,0,2,1,1,2,3,3,2,0,0,2,2,1,1,2,3,3,0,0,2,1,1,2,2,2,0,3,3,0))	;


	TYPE vec_array IS ARRAY (0 to 255, 0 to 15) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	TYPE vector_array IS ARRAY (0 to 7) OF vec_array;
-- constans used in P
	CONSTANT g512 : vector_array := (
	(
	(x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000"),
	(x"ef0b0270", x"3afd0000", x"5dae0000", x"69490000", x"9b0f3c06", x"4405b5f9", x"66140a51", x"924f5d0a", x"c96b0030", x"e7250000", x"2f840000", x"264f0000", x"08695bf9", x"6dfcf137", x"509f6984", x"9e69af68"),
	(x"c96b0030", x"e7250000", x"2f840000", x"264f0000", x"08695bf9", x"6dfcf137", x"509f6984", x"9e69af68", x"26600240", x"ddd80000", x"722a0000", x"4f060000", x"936667ff", x"29f944ce", x"368b63d5", x"0c26f262"),
	(x"26600240", x"ddd80000", x"722a0000", x"4f060000", x"936667ff", x"29f944ce", x"368b63d5", x"0c26f262", x"ef0b0270", x"3afd0000", x"5dae0000", x"69490000", x"9b0f3c06", x"4405b5f9", x"66140a51", x"924f5d0a"),
	(x"145a3c00", x"b9e90000", x"61270000", x"f1610000", x"ce613d6c", x"b0493d78", x"47a96720", x"e18e24c5", x"23671400", x"c8b90000", x"f4c70000", x"fb750000", x"73cd2465", x"f8a6a549", x"02c40a3f", x"dc24e61f"),
	(x"fb513e70", x"83140000", x"3c890000", x"98280000", x"556e016a", x"f44c8881", x"21bd6d71", x"73c179cf", x"ea0c1430", x"2f9c0000", x"db430000", x"dd3a0000", x"7ba47f9c", x"955a547e", x"525b63bb", x"424d4977"),
	(x"dd313c30", x"5ecc0000", x"4ea30000", x"d72e0000", x"c6086695", x"ddb5cc4f", x"17360ea4", x"7fe78bad", x"05071640", x"15610000", x"86ed0000", x"b4730000", x"e0ab439a", x"d15fe187", x"344f69ea", x"d002147d"),
	(x"323a3e40", x"64310000", x"130d0000", x"be670000", x"5d075a93", x"99b079b6", x"712204f5", x"eda8d6a7", x"cc6c1670", x"f2440000", x"a9690000", x"923c0000", x"e8c21863", x"bca310b0", x"64d0006e", x"4e6bbb15"),
	(x"23671400", x"c8b90000", x"f4c70000", x"fb750000", x"73cd2465", x"f8a6a549", x"02c40a3f", x"dc24e61f", x"373d2800", x"71500000", x"95e00000", x"0a140000", x"bdac1909", x"48ef9831", x"456d6d1f", x"3daac2da"),
	(x"cc6c1670", x"f2440000", x"a9690000", x"923c0000", x"e8c21863", x"bca310b0", x"64d0006e", x"4e6bbb15", x"fe562830", x"96750000", x"ba640000", x"2c5b0000", x"b5c542f0", x"25136906", x"15f2049b", x"a3c36db2"),
	(x"ea0c1430", x"2f9c0000", x"db430000", x"dd3a0000", x"7ba47f9c", x"955a547e", x"525b63bb", x"424d4977", x"115d2a40", x"ac880000", x"e7ca0000", x"45120000", x"2eca7ef6", x"6116dcff", x"73e60eca", x"318c30b8"),
	(x"05071640", x"15610000", x"86ed0000", x"b4730000", x"e0ab439a", x"d15fe187", x"344f69ea", x"d002147d", x"d8362a70", x"4bad0000", x"c84e0000", x"635d0000", x"26a3250f", x"0cea2dc8", x"2379674e", x"afe59fd0"),
	(x"373d2800", x"71500000", x"95e00000", x"0a140000", x"bdac1909", x"48ef9831", x"456d6d1f", x"3daac2da", x"145a3c00", x"b9e90000", x"61270000", x"f1610000", x"ce613d6c", x"b0493d78", x"47a96720", x"e18e24c5"),
	(x"d8362a70", x"4bad0000", x"c84e0000", x"635d0000", x"26a3250f", x"0cea2dc8", x"2379674e", x"afe59fd0", x"dd313c30", x"5ecc0000", x"4ea30000", x"d72e0000", x"c6086695", x"ddb5cc4f", x"17360ea4", x"7fe78bad"),
	(x"fe562830", x"96750000", x"ba640000", x"2c5b0000", x"b5c542f0", x"25136906", x"15f2049b", x"a3c36db2", x"323a3e40", x"64310000", x"130d0000", x"be670000", x"5d075a93", x"99b079b6", x"712204f5", x"eda8d6a7"),
	(x"115d2a40", x"ac880000", x"e7ca0000", x"45120000", x"2eca7ef6", x"6116dcff", x"73e60eca", x"318c30b8", x"fb513e70", x"83140000", x"3c890000", x"98280000", x"556e016a", x"f44c8881", x"21bd6d71", x"73c179cf"),
	(x"54285c00", x"eaed0000", x"c5d60000", x"a1c50000", x"b3a26770", x"94a5c4e1", x"6bb0419d", x"551b3782", x"9cbb1800", x"b0d30000", x"92510000", x"ed930000", x"593a4345", x"e114d5f4", x"430633da", x"78cace29"),
	(x"bb235e70", x"d0100000", x"98780000", x"c88c0000", x"28ad5b76", x"d0a07118", x"0da44bcc", x"c7546a88", x"55d01830", x"57f60000", x"bdd50000", x"cbdc0000", x"515318bc", x"8ce824c3", x"13995a5e", x"e6a36141"),
	(x"9d435c30", x"0dc80000", x"ea520000", x"878a0000", x"bbcb3c89", x"f95935d6", x"3b2f2819", x"cb7298ea", x"badb1a40", x"6d0b0000", x"e07b0000", x"a2950000", x"ca5c24ba", x"c8ed913a", x"758d500f", x"74ec3c4b"),
	(x"72485e40", x"37350000", x"b7fc0000", x"eec30000", x"20c4008f", x"bd5c802f", x"5d3b2248", x"593dc5e0", x"73b01a70", x"8a2e0000", x"cfff0000", x"84da0000", x"c2357f43", x"a511600d", x"2512398b", x"ea859323"),
	(x"40726000", x"53040000", x"a4f10000", x"50a40000", x"7dc35a1c", x"24ecf999", x"2c1926bd", x"b4951347", x"bfdc0c00", x"786a0000", x"66960000", x"16e60000", x"2af76720", x"19b270bd", x"41c239e5", x"a4ee2836"),
	(x"af796270", x"69f90000", x"f95f0000", x"39ed0000", x"e6cc661a", x"60e94c60", x"4a0d2cec", x"26da4e4d", x"76b70c30", x"9f4f0000", x"49120000", x"30a90000", x"229e3cd9", x"744e818a", x"115d5061", x"3a87875e"),
	(x"89196030", x"b4210000", x"8b750000", x"76eb0000", x"75aa01e5", x"491008ae", x"7c864f39", x"2afcbc2f", x"99bc0e40", x"a5b20000", x"14bc0000", x"59e00000", x"b99100df", x"304b3473", x"77495a30", x"a8c8da54"),
	(x"66126240", x"8edc0000", x"d6db0000", x"1fa20000", x"eea53de3", x"0d15bd57", x"1a924568", x"b8b3e125", x"50d70e70", x"42970000", x"3b380000", x"7faf0000", x"b1f85b26", x"5db7c544", x"27d633b4", x"36a1753c"),
	(x"774f4800", x"22540000", x"31110000", x"5ab00000", x"c06f4315", x"6c0361a8", x"69744ba2", x"893fd19d", x"ab863000", x"c1830000", x"07b10000", x"e7870000", x"e4965a4c", x"a9fb4dc5", x"066b5ec5", x"45600cf3"),
	(x"98444a70", x"18a90000", x"6cbf0000", x"33f90000", x"5b607f13", x"2806d451", x"0f6041f3", x"1b708c97", x"62ed3030", x"26a60000", x"28350000", x"c1c80000", x"ecff01b5", x"c407bcf2", x"56f43741", x"db09a39b"),
	(x"be244830", x"c5710000", x"1e950000", x"7cff0000", x"c80618ec", x"01ff909f", x"39eb2226", x"17567ef5", x"8de63240", x"1c5b0000", x"759b0000", x"a8810000", x"77f03db3", x"8002090b", x"30e03d10", x"4946fe91"),
	(x"512f4a40", x"ff8c0000", x"433b0000", x"15b60000", x"530924ea", x"45fa2566", x"5fff2877", x"851923ff", x"448d3270", x"fb7e0000", x"5a1f0000", x"8ece0000", x"7f99664a", x"edfef83c", x"607f5494", x"d72f51f9"),
	(x"63157400", x"9bbd0000", x"50360000", x"abd10000", x"0e0e7e79", x"dc4a5cd0", x"2edd2c82", x"68b1f558", x"88e12400", x"093a0000", x"f3760000", x"1cf20000", x"975b7e29", x"515de88c", x"04af54fa", x"9944eaec"),
	(x"8c1e7670", x"a1400000", x"0d980000", x"c2980000", x"9501427f", x"984fe929", x"48c926d3", x"fafea852", x"418a2430", x"ee1f0000", x"dcf20000", x"3abd0000", x"9f3225d0", x"3ca119bb", x"54303d7e", x"072d4584"),
	(x"aa7e7430", x"7c980000", x"7fb20000", x"8d9e0000", x"06672580", x"b1b6ade7", x"7e424506", x"f6d85a30", x"ae812640", x"d4e20000", x"815c0000", x"53f40000", x"043d19d6", x"78a4ac42", x"3224372f", x"9562188e"),
	(x"45757640", x"46650000", x"221c0000", x"e4d70000", x"9d681986", x"f5b3181e", x"18564f57", x"6497073a", x"67ea2670", x"33c70000", x"aed80000", x"75bb0000", x"0c54422f", x"15585d75", x"62bb5eab", x"0b0bb7e6"),
	(x"9cbb1800", x"b0d30000", x"92510000", x"ed930000", x"593a4345", x"e114d5f4", x"430633da", x"78cace29", x"c8934400", x"5a3e0000", x"57870000", x"4c560000", x"ea982435", x"75b11115", x"28b67247", x"2dd1f9ab"),
	(x"73b01a70", x"8a2e0000", x"cfff0000", x"84da0000", x"c2357f43", x"a511600d", x"2512398b", x"ea859323", x"01f84430", x"bd1b0000", x"78030000", x"6a190000", x"e2f17fcc", x"184de022", x"78291bc3", x"b3b856c3"),
	(x"55d01830", x"57f60000", x"bdd50000", x"cbdc0000", x"515318bc", x"8ce824c3", x"13995a5e", x"e6a36141", x"eef34640", x"87e60000", x"25ad0000", x"03500000", x"79fe43ca", x"5c4855db", x"1e3d1192", x"21f70bc9"),
	(x"badb1a40", x"6d0b0000", x"e07b0000", x"a2950000", x"ca5c24ba", x"c8ed913a", x"758d500f", x"74ec3c4b", x"27984670", x"60c30000", x"0a290000", x"251f0000", x"71971833", x"31b4a4ec", x"4ea27816", x"bf9ea4a1"),
	(x"88e12400", x"093a0000", x"f3760000", x"1cf20000", x"975b7e29", x"515de88c", x"04af54fa", x"9944eaec", x"ebf45000", x"92870000", x"a3400000", x"b7230000", x"99550050", x"8d17b45c", x"2a727878", x"f1f51fb4"),
	(x"67ea2670", x"33c70000", x"aed80000", x"75bb0000", x"0c54422f", x"15585d75", x"62bb5eab", x"0b0bb7e6", x"229f5030", x"75a20000", x"8cc40000", x"916c0000", x"913c5ba9", x"e0eb456b", x"7aed11fc", x"6f9cb0dc"),
	(x"418a2430", x"ee1f0000", x"dcf20000", x"3abd0000", x"9f3225d0", x"3ca119bb", x"54303d7e", x"072d4584", x"cd945240", x"4f5f0000", x"d16a0000", x"f8250000", x"0a3367af", x"a4eef092", x"1cf91bad", x"fdd3edd6"),
	(x"ae812640", x"d4e20000", x"815c0000", x"53f40000", x"043d19d6", x"78a4ac42", x"3224372f", x"9562188e", x"04ff5270", x"a87a0000", x"feee0000", x"de6a0000", x"025a3c56", x"c91201a5", x"4c667229", x"63ba42be"),
	(x"bfdc0c00", x"786a0000", x"66960000", x"16e60000", x"2af76720", x"19b270bd", x"41c239e5", x"a4ee2836", x"ffae6c00", x"2b6e0000", x"c2670000", x"46420000", x"57343d3c", x"3d5e8924", x"6ddb1f58", x"107b3b71"),
	(x"50d70e70", x"42970000", x"3b380000", x"7faf0000", x"b1f85b26", x"5db7c544", x"27d633b4", x"36a1753c", x"36c56c30", x"cc4b0000", x"ede30000", x"600d0000", x"5f5d66c5", x"50a27813", x"3d4476dc", x"8e129419"),
	(x"76b70c30", x"9f4f0000", x"49120000", x"30a90000", x"229e3cd9", x"744e818a", x"115d5061", x"3a87875e", x"d9ce6e40", x"f6b60000", x"b04d0000", x"09440000", x"c4525ac3", x"14a7cdea", x"5b507c8d", x"1c5dc913"),
	(x"99bc0e40", x"a5b20000", x"14bc0000", x"59e00000", x"b99100df", x"304b3473", x"77495a30", x"a8c8da54", x"10a56e70", x"11930000", x"9fc90000", x"2f0b0000", x"cc3b013a", x"795b3cdd", x"0bcf1509", x"8234667b"),
	(x"ab863000", x"c1830000", x"07b10000", x"e7870000", x"e4965a4c", x"a9fb4dc5", x"066b5ec5", x"45600cf3", x"dcc97800", x"e3d70000", x"36a00000", x"bd370000", x"24f91959", x"c5f82c6d", x"6f1f1567", x"cc5fdd6e"),
	(x"448d3270", x"fb7e0000", x"5a1f0000", x"8ece0000", x"7f99664a", x"edfef83c", x"607f5494", x"d72f51f9", x"15a27830", x"04f20000", x"19240000", x"9b780000", x"2c9042a0", x"a804dd5a", x"3f807ce3", x"52367206"),
	(x"62ed3030", x"26a60000", x"28350000", x"c1c80000", x"ecff01b5", x"c407bcf2", x"56f43741", x"db09a39b", x"faa97a40", x"3e0f0000", x"448a0000", x"f2310000", x"b79f7ea6", x"ec0168a3", x"599476b2", x"c0792f0c"),
	(x"8de63240", x"1c5b0000", x"759b0000", x"a8810000", x"77f03db3", x"8002090b", x"30e03d10", x"4946fe91", x"33c27a70", x"d92a0000", x"6b0e0000", x"d47e0000", x"bff6255f", x"81fd9994", x"090b1f36", x"5e108064"),
	(x"c8934400", x"5a3e0000", x"57870000", x"4c560000", x"ea982435", x"75b11115", x"28b67247", x"2dd1f9ab", x"54285c00", x"eaed0000", x"c5d60000", x"a1c50000", x"b3a26770", x"94a5c4e1", x"6bb0419d", x"551b3782"),
	(x"27984670", x"60c30000", x"0a290000", x"251f0000", x"71971833", x"31b4a4ec", x"4ea27816", x"bf9ea4a1", x"9d435c30", x"0dc80000", x"ea520000", x"878a0000", x"bbcb3c89", x"f95935d6", x"3b2f2819", x"cb7298ea"),
	(x"01f84430", x"bd1b0000", x"78030000", x"6a190000", x"e2f17fcc", x"184de022", x"78291bc3", x"b3b856c3", x"72485e40", x"37350000", x"b7fc0000", x"eec30000", x"20c4008f", x"bd5c802f", x"5d3b2248", x"593dc5e0"),
	(x"eef34640", x"87e60000", x"25ad0000", x"03500000", x"79fe43ca", x"5c4855db", x"1e3d1192", x"21f70bc9", x"bb235e70", x"d0100000", x"98780000", x"c88c0000", x"28ad5b76", x"d0a07118", x"0da44bcc", x"c7546a88"),
	(x"dcc97800", x"e3d70000", x"36a00000", x"bd370000", x"24f91959", x"c5f82c6d", x"6f1f1567", x"cc5fdd6e", x"774f4800", x"22540000", x"31110000", x"5ab00000", x"c06f4315", x"6c0361a8", x"69744ba2", x"893fd19d"),
	(x"33c27a70", x"d92a0000", x"6b0e0000", x"d47e0000", x"bff6255f", x"81fd9994", x"090b1f36", x"5e108064", x"be244830", x"c5710000", x"1e950000", x"7cff0000", x"c80618ec", x"01ff909f", x"39eb2226", x"17567ef5"),
	(x"15a27830", x"04f20000", x"19240000", x"9b780000", x"2c9042a0", x"a804dd5a", x"3f807ce3", x"52367206", x"512f4a40", x"ff8c0000", x"433b0000", x"15b60000", x"530924ea", x"45fa2566", x"5fff2877", x"851923ff"),
	(x"faa97a40", x"3e0f0000", x"448a0000", x"f2310000", x"b79f7ea6", x"ec0168a3", x"599476b2", x"c0792f0c", x"98444a70", x"18a90000", x"6cbf0000", x"33f90000", x"5b607f13", x"2806d451", x"0f6041f3", x"1b708c97"),
	(x"ebf45000", x"92870000", x"a3400000", x"b7230000", x"99550050", x"8d17b45c", x"2a727878", x"f1f51fb4", x"63157400", x"9bbd0000", x"50360000", x"abd10000", x"0e0e7e79", x"dc4a5cd0", x"2edd2c82", x"68b1f558"),
	(x"04ff5270", x"a87a0000", x"feee0000", x"de6a0000", x"025a3c56", x"c91201a5", x"4c667229", x"63ba42be", x"aa7e7430", x"7c980000", x"7fb20000", x"8d9e0000", x"06672580", x"b1b6ade7", x"7e424506", x"f6d85a30"),
	(x"229f5030", x"75a20000", x"8cc40000", x"916c0000", x"913c5ba9", x"e0eb456b", x"7aed11fc", x"6f9cb0dc", x"45757640", x"46650000", x"221c0000", x"e4d70000", x"9d681986", x"f5b3181e", x"18564f57", x"6497073a"),
	(x"cd945240", x"4f5f0000", x"d16a0000", x"f8250000", x"0a3367af", x"a4eef092", x"1cf91bad", x"fdd3edd6", x"8c1e7670", x"a1400000", x"0d980000", x"c2980000", x"9501427f", x"984fe929", x"48c926d3", x"fafea852"),
	(x"ffae6c00", x"2b6e0000", x"c2670000", x"46420000", x"57343d3c", x"3d5e8924", x"6ddb1f58", x"107b3b71", x"40726000", x"53040000", x"a4f10000", x"50a40000", x"7dc35a1c", x"24ecf999", x"2c1926bd", x"b4951347"),
	(x"10a56e70", x"11930000", x"9fc90000", x"2f0b0000", x"cc3b013a", x"795b3cdd", x"0bcf1509", x"8234667b", x"89196030", x"b4210000", x"8b750000", x"76eb0000", x"75aa01e5", x"491008ae", x"7c864f39", x"2afcbc2f"),
	(x"36c56c30", x"cc4b0000", x"ede30000", x"600d0000", x"5f5d66c5", x"50a27813", x"3d4476dc", x"8e129419", x"66126240", x"8edc0000", x"d6db0000", x"1fa20000", x"eea53de3", x"0d15bd57", x"1a924568", x"b8b3e125"),
	(x"d9ce6e40", x"f6b60000", x"b04d0000", x"09440000", x"c4525ac3", x"14a7cdea", x"5b507c8d", x"1c5dc913", x"af796270", x"69f90000", x"f95f0000", x"39ed0000", x"e6cc661a", x"60e94c60", x"4a0d2cec", x"26da4e4d"),
	(x"29449c00", x"64e70000", x"f24b0000", x"c2f30000", x"0ede4e8f", x"56c23745", x"f3e04259", x"8d0d9ec4", x"466d0c00", x"08620000", x"dd5d0000", x"badd0000", x"6a927942", x"441f2b93", x"218ace6f", x"bf2c0be2"),
	(x"c64f9e70", x"5e1a0000", x"afe50000", x"abba0000", x"95d17289", x"12c782bc", x"95f44808", x"1f42c3ce", x"8f060c30", x"ef470000", x"f2d90000", x"9c920000", x"62fb22bb", x"29e3daa4", x"7115a7eb", x"2145a48a"),
	(x"e02f9c30", x"83c20000", x"ddcf0000", x"e4bc0000", x"06b71576", x"3b3ec672", x"a37f2bdd", x"136431ac", x"600d0e40", x"d5ba0000", x"af770000", x"f5db0000", x"f9f41ebd", x"6de66f5d", x"1701adba", x"b30af980"),
	(x"0f249e40", x"b93f0000", x"80610000", x"8df50000", x"9db82970", x"7f3b738b", x"c56b218c", x"812b6ca6", x"a9660e70", x"329f0000", x"80f30000", x"d3940000", x"f19d4544", x"001a9e6a", x"479ec43e", x"2d6356e8"),
	(x"3d1ea000", x"dd0e0000", x"936c0000", x"33920000", x"c0bf73e3", x"e68b0a3d", x"b4492579", x"6c83ba01", x"650a1800", x"c0db0000", x"299a0000", x"41a80000", x"195f5d27", x"bcb98eda", x"234ec450", x"6308edfd"),
	(x"d215a270", x"e7f30000", x"cec20000", x"5adb0000", x"5bb04fe5", x"a28ebfc4", x"d25d2f28", x"fecce70b", x"ac611830", x"27fe0000", x"061e0000", x"67e70000", x"113606de", x"d1457fed", x"73d1add4", x"fd614295"),
	(x"f475a030", x"3a2b0000", x"bce80000", x"15dd0000", x"c8d6281a", x"8b77fb0a", x"e4d64cfd", x"f2ea1569", x"436a1a40", x"1d030000", x"5bb00000", x"0eae0000", x"8a393ad8", x"9540ca14", x"15c5a785", x"6f2e1f9f"),
	(x"1b7ea240", x"00d60000", x"e1460000", x"7c940000", x"53d9141c", x"cf724ef3", x"82c246ac", x"60a54863", x"8a011a70", x"fa260000", x"74340000", x"28e10000", x"82506121", x"f8bc3b23", x"455ace01", x"f147b0f7"),
	(x"0a238800", x"ac5e0000", x"068c0000", x"39860000", x"7d136aea", x"ae64920c", x"f1244866", x"512978db", x"71502400", x"79320000", x"48bd0000", x"b0c90000", x"d73e604b", x"0cf0b3a2", x"64e7a370", x"8286c938"),
	(x"e5288a70", x"96a30000", x"5b220000", x"50cf0000", x"e61c56ec", x"ea6127f5", x"97304237", x"c36625d1", x"b83b2430", x"9e170000", x"67390000", x"96860000", x"df573bb2", x"610c4295", x"3478caf4", x"1cef6650"),
	(x"c3488830", x"4b7b0000", x"29080000", x"1fc90000", x"757a3113", x"c398633b", x"a1bb21e2", x"cf40d7b3", x"57302640", x"a4ea0000", x"3a970000", x"ffcf0000", x"445807b4", x"2509f76c", x"526cc0a5", x"8ea03b5a"),
	(x"2c438a40", x"71860000", x"74a60000", x"76800000", x"ee750d15", x"879dd6c2", x"c7af2bb3", x"5d0f8ab9", x"9e5b2670", x"43cf0000", x"15130000", x"d9800000", x"4c315c4d", x"48f5065b", x"02f3a921", x"10c99432"),
	(x"1e79b400", x"15b70000", x"67ab0000", x"c8e70000", x"b3725786", x"1e2daf74", x"b68d2f46", x"b0a75c1e", x"52373000", x"b18b0000", x"bc7a0000", x"4bbc0000", x"a4f3442e", x"f45616eb", x"6623a94f", x"5ea22f27"),
	(x"f172b670", x"2f4a0000", x"3a050000", x"a1ae0000", x"287d6b80", x"5a281a8d", x"d0992517", x"22e80114", x"9b5c3030", x"56ae0000", x"93fe0000", x"6df30000", x"ac9a1fd7", x"99aae7dc", x"36bcc0cb", x"c0cb804f"),
	(x"d712b430", x"f2920000", x"482f0000", x"eea80000", x"bb1b0c7f", x"73d15e43", x"e61246c2", x"2ecef376", x"74573240", x"6c530000", x"ce500000", x"04ba0000", x"379523d1", x"ddaf5225", x"50a8ca9a", x"5284dd45"),
	(x"3819b640", x"c86f0000", x"15810000", x"87e10000", x"20143079", x"37d4ebba", x"80064c93", x"bc81ae7c", x"bd3c3270", x"8b760000", x"e1d40000", x"22f50000", x"3ffc7828", x"b053a312", x"0037a31e", x"cced722d"),
	(x"7d6cc000", x"8e0a0000", x"379d0000", x"63360000", x"bd7c29ff", x"c267f3a4", x"985003c4", x"d816a946", x"dad61400", x"b8b10000", x"4f0c0000", x"574e0000", x"33a83a07", x"a50bfe67", x"628cfdb5", x"c7e6c5cb"),
	(x"9267c270", x"b4f70000", x"6a330000", x"0a7f0000", x"267315f9", x"8662465d", x"fe440995", x"4a59f44c", x"13bd1430", x"5f940000", x"60880000", x"71010000", x"3bc161fe", x"c8f70f50", x"32139431", x"598f6aa3"),
	(x"b407c030", x"692f0000", x"18190000", x"45790000", x"b5157206", x"af9b0293", x"c8cf6a40", x"467f062e", x"fcb61640", x"65690000", x"3d260000", x"18480000", x"a0ce5df8", x"8cf2baa9", x"54079e60", x"cbc037a9"),
	(x"5b0cc240", x"53d20000", x"45b70000", x"2c300000", x"2e1a4e00", x"eb9eb76a", x"aedb6011", x"d4305b24", x"35dd1670", x"824c0000", x"12a20000", x"3e070000", x"a8a70601", x"e10e4b9e", x"0498f7e4", x"55a998c1"),
	(x"6936fc00", x"37e30000", x"56ba0000", x"92570000", x"731d1493", x"722ecedc", x"dff964e4", x"39988d83", x"f9b10000", x"70080000", x"bbcb0000", x"ac3b0000", x"40651e62", x"5dad5b2e", x"6048f78a", x"1bc223d4"),
	(x"863dfe70", x"0d1e0000", x"0b140000", x"fb1e0000", x"e8122895", x"362b7b25", x"b9ed6eb5", x"abd7d089", x"30da0030", x"972d0000", x"944f0000", x"8a740000", x"480c459b", x"3051aa19", x"30d79e0e", x"85ab8cbc"),
	(x"a05dfc30", x"d0c60000", x"793e0000", x"b4180000", x"7b744f6a", x"1fd23feb", x"8f660d60", x"a7f122eb", x"dfd10240", x"add00000", x"c9e10000", x"e33d0000", x"d303799d", x"74541fe0", x"56c3945f", x"17e4d1b6"),
	(x"4f56fe40", x"ea3b0000", x"24900000", x"dd510000", x"e07b736c", x"5bd78a12", x"e9720731", x"35be7fe1", x"16ba0270", x"4af50000", x"e6650000", x"c5720000", x"db6a2264", x"19a8eed7", x"065cfddb", x"898d7ede"),
	(x"5e0bd400", x"46b30000", x"c35a0000", x"98430000", x"ceb10d9a", x"3ac156ed", x"9a9409fb", x"04324f59", x"edeb3c00", x"c9e10000", x"daec0000", x"5d5a0000", x"8e04230e", x"ede46656", x"27e190aa", x"fa4c0711"),
	(x"b100d670", x"7c4e0000", x"9ef40000", x"f10a0000", x"55be319c", x"7ec4e314", x"fc8003aa", x"967d1253", x"24803c30", x"2ec40000", x"f5680000", x"7b150000", x"866d78f7", x"80189761", x"777ef92e", x"6425a879"),
	(x"9760d430", x"a1960000", x"ecde0000", x"be0c0000", x"c6d85663", x"573da7da", x"ca0b607f", x"9a5be031", x"cb8b3e40", x"14390000", x"a8c60000", x"125c0000", x"1d6244f1", x"c41d2298", x"116af37f", x"f66af573"),
	(x"786bd640", x"9b6b0000", x"b1700000", x"d7450000", x"5dd76a65", x"13381223", x"ac1f6a2e", x"0814bd3b", x"02e03e70", x"f31c0000", x"87420000", x"34130000", x"150b1f08", x"a9e1d3af", x"41f59afb", x"68035a1b"),
	(x"4a51e800", x"ff5a0000", x"a27d0000", x"69220000", x"00d030f6", x"8a886b95", x"dd3d6edb", x"e5bc6b9c", x"ce8c2800", x"01580000", x"2e2b0000", x"a62f0000", x"fdc9076b", x"1542c31f", x"25259a95", x"2668e10e"),
	(x"a55aea70", x"c5a70000", x"ffd30000", x"006b0000", x"9bdf0cf0", x"ce8dde6c", x"bb29648a", x"77f33696", x"07e72830", x"e67d0000", x"01af0000", x"80600000", x"f5a05c92", x"78be3228", x"75baf311", x"b8014e66"),
	(x"833ae830", x"187f0000", x"8df90000", x"4f6d0000", x"08b96b0f", x"e7749aa2", x"8da2075f", x"7bd5c4f4", x"e8ec2a40", x"dc800000", x"5c010000", x"e9290000", x"6eaf6094", x"3cbb87d1", x"13aef940", x"2a4e136c"),
	(x"6c31ea40", x"22820000", x"d0570000", x"26240000", x"93b65709", x"a3712f5b", x"ebb60d0e", x"e99a99fe", x"21872a70", x"3ba50000", x"73850000", x"cf660000", x"66c63b6d", x"514776e6", x"433190c4", x"b427bc04"),
	(x"b5ff8400", x"d4340000", x"601a0000", x"2f600000", x"57e40dca", x"b7d6e2b1", x"b0e67183", x"f5c750ed", x"8efe4800", x"525c0000", x"8ada0000", x"f68b0000", x"800a5d77", x"31ae3a86", x"093cbc28", x"92fdf249"),
	(x"5af48670", x"eec90000", x"3db40000", x"46290000", x"cceb31cc", x"f3d35748", x"d6f27bd2", x"67880de7", x"47954830", x"b5790000", x"a55e0000", x"d0c40000", x"8863068e", x"5c52cbb1", x"59a3d5ac", x"0c945d21"),
	(x"7c948430", x"33110000", x"4f9e0000", x"092f0000", x"5f8d5633", x"da2a1386", x"e0791807", x"6baeff85", x"a89e4a40", x"8f840000", x"f8f00000", x"b98d0000", x"136c3a88", x"18577e48", x"3fb7dffd", x"9edb002b"),
	(x"939f8640", x"09ec0000", x"12300000", x"60660000", x"c4826a35", x"9e2fa67f", x"866d1256", x"f9e1a28f", x"61f54a70", x"68a10000", x"d7740000", x"9fc20000", x"1b056171", x"75ab8f7f", x"6f28b679", x"00b2af43"),
	(x"a1a5b800", x"6ddd0000", x"013d0000", x"de010000", x"998530a6", x"079fdfc9", x"f74f16a3", x"14497428", x"ad995c00", x"9ae50000", x"7e1d0000", x"0dfe0000", x"f3c77912", x"c9089fcf", x"0bf8b617", x"4ed91456"),
	(x"4eaeba70", x"57200000", x"5c930000", x"b7480000", x"028a0ca0", x"439a6a30", x"915b1cf2", x"86062922", x"64f25c30", x"7dc00000", x"51990000", x"2bb10000", x"fbae22eb", x"a4f46ef8", x"5b67df93", x"d0b0bb3e"),
	(x"68ceb830", x"8af80000", x"2eb90000", x"f84e0000", x"91ec6b5f", x"6a632efe", x"a7d07f27", x"8a20db40", x"8bf95e40", x"473d0000", x"0c370000", x"42f80000", x"60a11eed", x"e0f1db01", x"3d73d5c2", x"42ffe634"),
	(x"87c5ba40", x"b0050000", x"73170000", x"91070000", x"0ae35759", x"2e669b07", x"c1c47576", x"186f864a", x"42925e70", x"a0180000", x"23b30000", x"64b70000", x"68c84514", x"8d0d2a36", x"6decbc46", x"dc96495c"),
	(x"96989000", x"1c8d0000", x"94dd0000", x"d4150000", x"242929af", x"4f7047f8", x"b2227bbc", x"29e3b6f2", x"b9c36000", x"230c0000", x"1f3a0000", x"fc9f0000", x"3da6447e", x"7941a2b7", x"4c51d137", x"af573093"),
	(x"79939270", x"26700000", x"c9730000", x"bd5c0000", x"bf2615a9", x"0b75f201", x"d43671ed", x"bbacebf8", x"70a86030", x"c4290000", x"30be0000", x"dad00000", x"35cf1f87", x"14bd5380", x"1cceb8b3", x"313e9ffb"),
	(x"5ff39030", x"fba80000", x"bb590000", x"f25a0000", x"2c407256", x"228cb6cf", x"e2bd1238", x"b78a199a", x"9fa36240", x"fed40000", x"6d100000", x"b3990000", x"aec02381", x"50b8e679", x"7adab2e2", x"a371c2f1"),
	(x"b0f89240", x"c1550000", x"e6f70000", x"9b130000", x"b74f4e50", x"66890336", x"84a91869", x"25c54490", x"56c86270", x"19f10000", x"42940000", x"95d60000", x"a6a97878", x"3d44174e", x"2a45db66", x"3d186d99"),
	(x"82c2ac00", x"a5640000", x"f5fa0000", x"25740000", x"ea4814c3", x"ff397a80", x"f58b1c9c", x"c86d9237", x"9aa47400", x"ebb50000", x"ebfd0000", x"07ea0000", x"4e6b601b", x"81e707fe", x"4e95db08", x"7373d68c"),
	(x"6dc9ae70", x"9f990000", x"a8540000", x"4c3d0000", x"714728c5", x"bb3ccf79", x"939f16cd", x"5a22cf3d", x"53cf7430", x"0c900000", x"c4790000", x"21a50000", x"46023be2", x"ec1bf6c9", x"1e0ab28c", x"ed1a79e4"),
	(x"4ba9ac30", x"42410000", x"da7e0000", x"033b0000", x"e2214f3a", x"92c58bb7", x"a5147518", x"56043d5f", x"bcc47640", x"366d0000", x"99d70000", x"48ec0000", x"dd0d07e4", x"a81e4330", x"781eb8dd", x"7f5524ee"),
	(x"a4a2ae40", x"78bc0000", x"87d00000", x"6a720000", x"792e733c", x"d6c03e4e", x"c3007f49", x"c44b6055", x"75af7670", x"d1480000", x"b6530000", x"6ea30000", x"d5645c1d", x"c5e2b207", x"2881d159", x"e13c8b86"),
	(x"e1d7d800", x"3ed90000", x"a5cc0000", x"8ea50000", x"e4466aba", x"23732650", x"db56301e", x"a0dc676f", x"12455000", x"e28f0000", x"188b0000", x"1b180000", x"d9301e32", x"d0baef72", x"4a3a8ff2", x"ea373c60"),
	(x"0edcda70", x"04240000", x"f8620000", x"e7ec0000", x"7f4956bc", x"677693a9", x"bd423a4f", x"32933a65", x"db2e5030", x"05aa0000", x"370f0000", x"3d570000", x"d15945cb", x"bd461e45", x"1aa5e676", x"745e9308"),
	(x"28bcd830", x"d9fc0000", x"8a480000", x"a8ea0000", x"ec2f3143", x"4e8fd767", x"8bc9599a", x"3eb5c807", x"34255240", x"3f570000", x"6aa10000", x"541e0000", x"4a5679cd", x"f943abbc", x"7cb1ec27", x"e611ce02"),
	(x"c7b7da40", x"e3010000", x"d7e60000", x"c1a30000", x"77200d45", x"0a8a629e", x"eddd53cb", x"acfa950d", x"fd4e5270", x"d8720000", x"45250000", x"72510000", x"423f2234", x"94bf5a8b", x"2c2e85a3", x"7878616a"),
	(x"f58de400", x"87300000", x"c4eb0000", x"7fc40000", x"2a2757d6", x"933a1b28", x"9cff573e", x"415243aa", x"31224400", x"2a360000", x"ec4c0000", x"e06d0000", x"aafd3a57", x"281c4a3b", x"48fe85cd", x"3613da7f"),
	(x"1a86e670", x"bdcd0000", x"99450000", x"168d0000", x"b1286bd0", x"d73faed1", x"faeb5d6f", x"d31d1ea0", x"f8494430", x"cd130000", x"c3c80000", x"c6220000", x"a29461ae", x"45e0bb0c", x"1861ec49", x"a87a7517"),
	(x"3ce6e430", x"60150000", x"eb6f0000", x"598b0000", x"224e0c2f", x"fec6ea1f", x"cc603eba", x"df3becc2", x"17424640", x"f7ee0000", x"9e660000", x"af6b0000", x"399b5da8", x"01e50ef5", x"7e75e618", x"3a35281d"),
	(x"d3ede640", x"5ae80000", x"b6c10000", x"30c20000", x"b9413029", x"bac35fe6", x"aa7434eb", x"4d74b1c8", x"de294670", x"10cb0000", x"b1e20000", x"89240000", x"31f20651", x"6c19ffc2", x"2eea8f9c", x"a45c8775"),
	(x"c2b0cc00", x"f6600000", x"510b0000", x"75d00000", x"978b4edf", x"dbd58319", x"d9923a21", x"7cf88170", x"25787800", x"93df0000", x"8d6b0000", x"110c0000", x"649c073b", x"98557743", x"0f57e2ed", x"d79dfeba"),
	(x"2dbbce70", x"cc9d0000", x"0ca50000", x"1c990000", x"0c8472d9", x"9fd036e0", x"bf863070", x"eeb7dc7a", x"ec137830", x"74fa0000", x"a2ef0000", x"37430000", x"6cf55cc2", x"f5a98674", x"5fc88b69", x"49f451d2"),
	(x"0bdbcc30", x"11450000", x"7e8f0000", x"539f0000", x"9fe21526", x"b629722e", x"890d53a5", x"e2912e18", x"03187a40", x"4e070000", x"ff410000", x"5e0a0000", x"f7fa60c4", x"b1ac338d", x"39dc8138", x"dbbb0cd8"),
	(x"e4d0ce40", x"2bb80000", x"23210000", x"3ad60000", x"04ed2920", x"f22cc7d7", x"ef1959f4", x"70de7312", x"ca737a70", x"a9220000", x"d0c50000", x"78450000", x"ff933b3d", x"dc50c2ba", x"6943e8bc", x"45d2a3b0"),
	(x"d6eaf000", x"4f890000", x"302c0000", x"84b10000", x"59ea73b3", x"6b9cbe61", x"9e3b5d01", x"9d76a5b5", x"061f6c00", x"5b660000", x"79ac0000", x"ea790000", x"1751235e", x"60f3d20a", x"0d93e8d2", x"0bb918a5"),
	(x"39e1f270", x"75740000", x"6d820000", x"edf80000", x"c2e54fb5", x"2f990b98", x"f82f5750", x"0f39f8bf", x"cf746c30", x"bc430000", x"56280000", x"cc360000", x"1f3878a7", x"0d0f233d", x"5d0c8156", x"95d0b7cd"),
	(x"1f81f030", x"a8ac0000", x"1fa80000", x"a2fe0000", x"5183284a", x"06604f56", x"cea43485", x"031f0add", x"207f6e40", x"86be0000", x"0b860000", x"a57f0000", x"843744a1", x"490a96c4", x"3b188b07", x"079feac7"),
	(x"f08af240", x"92510000", x"42060000", x"cbb70000", x"ca8c144c", x"4265faaf", x"a8b03ed4", x"915057d7", x"e9146e70", x"619b0000", x"24020000", x"83300000", x"8c5e1f58", x"24f667f3", x"6b87e283", x"99f645af"),
	(x"466d0c00", x"08620000", x"dd5d0000", x"badd0000", x"6a927942", x"441f2b93", x"218ace6f", x"bf2c0be2", x"6f299000", x"6c850000", x"2f160000", x"782e0000", x"644c37cd", x"12dd1cd6", x"d26a8c36", x"32219526"),
	(x"a9660e70", x"329f0000", x"80f30000", x"d3940000", x"f19d4544", x"001a9e6a", x"479ec43e", x"2d6356e8", x"a6429030", x"8ba00000", x"00920000", x"5e610000", x"6c256c34", x"7f21ede1", x"82f5e5b2", x"ac483a4e"),
	(x"8f060c30", x"ef470000", x"f2d90000", x"9c920000", x"62fb22bb", x"29e3daa4", x"7115a7eb", x"2145a48a", x"49499240", x"b15d0000", x"5d3c0000", x"37280000", x"f72a5032", x"3b245818", x"e4e1efe3", x"3e076744"),
	(x"600d0e40", x"d5ba0000", x"af770000", x"f5db0000", x"f9f41ebd", x"6de66f5d", x"1701adba", x"b30af980", x"80229270", x"56780000", x"72b80000", x"11670000", x"ff430bcb", x"56d8a92f", x"b47e8667", x"a06ec82c"),
	(x"52373000", x"b18b0000", x"bc7a0000", x"4bbc0000", x"a4f3442e", x"f45616eb", x"6623a94f", x"5ea22f27", x"4c4e8400", x"a43c0000", x"dbd10000", x"835b0000", x"178113a8", x"ea7bb99f", x"d0ae8609", x"ee057339"),
	(x"bd3c3270", x"8b760000", x"e1d40000", x"22f50000", x"3ffc7828", x"b053a312", x"0037a31e", x"cced722d", x"85258430", x"43190000", x"f4550000", x"a5140000", x"1fe84851", x"878748a8", x"8031ef8d", x"706cdc51"),
	(x"9b5c3030", x"56ae0000", x"93fe0000", x"6df30000", x"ac9a1fd7", x"99aae7dc", x"36bcc0cb", x"c0cb804f", x"6a2e8640", x"79e40000", x"a9fb0000", x"cc5d0000", x"84e77457", x"c382fd51", x"e625e5dc", x"e223815b"),
	(x"74573240", x"6c530000", x"ce500000", x"04ba0000", x"379523d1", x"ddaf5225", x"50a8ca9a", x"5284dd45", x"a3458670", x"9ec10000", x"867f0000", x"ea120000", x"8c8e2fae", x"ae7e0c66", x"b6ba8c58", x"7c4a2e33"),
	(x"650a1800", x"c0db0000", x"299a0000", x"41a80000", x"195f5d27", x"bcb98eda", x"234ec450", x"6308edfd", x"5814b800", x"1dd50000", x"baf60000", x"723a0000", x"d9e02ec4", x"5a3284e7", x"9707e129", x"0f8b57fc"),
	(x"8a011a70", x"fa260000", x"74340000", x"28e10000", x"82506121", x"f8bc3b23", x"455ace01", x"f147b0f7", x"917fb830", x"faf00000", x"95720000", x"54750000", x"d189753d", x"37ce75d0", x"c79888ad", x"91e2f894"),
	(x"ac611830", x"27fe0000", x"061e0000", x"67e70000", x"113606de", x"d1457fed", x"73d1add4", x"fd614295", x"7e74ba40", x"c00d0000", x"c8dc0000", x"3d3c0000", x"4a86493b", x"73cbc029", x"a18c82fc", x"03ada59e"),
	(x"436a1a40", x"1d030000", x"5bb00000", x"0eae0000", x"8a393ad8", x"9540ca14", x"15c5a785", x"6f2e1f9f", x"b71fba70", x"27280000", x"e7580000", x"1b730000", x"42ef12c2", x"1e37311e", x"f113eb78", x"9dc40af6"),
	(x"71502400", x"79320000", x"48bd0000", x"b0c90000", x"d73e604b", x"0cf0b3a2", x"64e7a370", x"8286c938", x"7b73ac00", x"d56c0000", x"4e310000", x"894f0000", x"aa2d0aa1", x"a29421ae", x"95c3eb16", x"d3afb1e3"),
	(x"9e5b2670", x"43cf0000", x"15130000", x"d9800000", x"4c315c4d", x"48f5065b", x"02f3a921", x"10c99432", x"b218ac30", x"32490000", x"61b50000", x"af000000", x"a2445158", x"cf68d099", x"c55c8292", x"4dc61e8b"),
	(x"b83b2430", x"9e170000", x"67390000", x"96860000", x"df573bb2", x"610c4295", x"3478caf4", x"1cef6650", x"5d13ae40", x"08b40000", x"3c1b0000", x"c6490000", x"394b6d5e", x"8b6d6560", x"a34888c3", x"df894381"),
	(x"57302640", x"a4ea0000", x"3a970000", x"ffcf0000", x"445807b4", x"2509f76c", x"526cc0a5", x"8ea03b5a", x"9478ae70", x"ef910000", x"139f0000", x"e0060000", x"312236a7", x"e6919457", x"f3d7e147", x"41e0ece9"),
	(x"12455000", x"e28f0000", x"188b0000", x"1b180000", x"d9301e32", x"d0baef72", x"4a3a8ff2", x"ea373c60", x"f3928800", x"dc560000", x"bd470000", x"95bd0000", x"3d767488", x"f3c9c922", x"916cbfec", x"4aeb5b0f"),
	(x"fd4e5270", x"d8720000", x"45250000", x"72510000", x"423f2234", x"94bf5a8b", x"2c2e85a3", x"7878616a", x"3af98830", x"3b730000", x"92c30000", x"b3f20000", x"351f2f71", x"9e353815", x"c1f3d668", x"d482f467"),
	(x"db2e5030", x"05aa0000", x"370f0000", x"3d570000", x"d15945cb", x"bd461e45", x"1aa5e676", x"745e9308", x"d5f28a40", x"018e0000", x"cf6d0000", x"dabb0000", x"ae101377", x"da308dec", x"a7e7dc39", x"46cda96d"),
	(x"34255240", x"3f570000", x"6aa10000", x"541e0000", x"4a5679cd", x"f943abbc", x"7cb1ec27", x"e611ce02", x"1c998a70", x"e6ab0000", x"e0e90000", x"fcf40000", x"a679488e", x"b7cc7cdb", x"f778b5bd", x"d8a40605"),
	(x"061f6c00", x"5b660000", x"79ac0000", x"ea790000", x"1751235e", x"60f3d20a", x"0d93e8d2", x"0bb918a5", x"d0f59c00", x"14ef0000", x"49800000", x"6ec80000", x"4ebb50ed", x"0b6f6c6b", x"93a8b5d3", x"96cfbd10"),
	(x"e9146e70", x"619b0000", x"24020000", x"83300000", x"8c5e1f58", x"24f667f3", x"6b87e283", x"99f645af", x"199e9c30", x"f3ca0000", x"66040000", x"48870000", x"46d20b14", x"66939d5c", x"c337dc57", x"08a61278"),
	(x"cf746c30", x"bc430000", x"56280000", x"cc360000", x"1f3878a7", x"0d0f233d", x"5d0c8156", x"95d0b7cd", x"f6959e40", x"c9370000", x"3baa0000", x"21ce0000", x"dddd3712", x"229628a5", x"a523d606", x"9ae94f72"),
	(x"207f6e40", x"86be0000", x"0b860000", x"a57f0000", x"843744a1", x"490a96c4", x"3b188b07", x"079feac7", x"3ffe9e70", x"2e120000", x"142e0000", x"07810000", x"d5b46ceb", x"4f6ad992", x"f5bcbf82", x"0480e01a"),
	(x"31224400", x"2a360000", x"ec4c0000", x"e06d0000", x"aafd3a57", x"281c4a3b", x"48fe85cd", x"3613da7f", x"c4afa000", x"ad060000", x"28a70000", x"9fa90000", x"80da6d81", x"bb265113", x"d401d2f3", x"774199d5"),
	(x"de294670", x"10cb0000", x"b1e20000", x"89240000", x"31f20651", x"6c19ffc2", x"2eea8f9c", x"a45c8775", x"0dc4a030", x"4a230000", x"07230000", x"b9e60000", x"88b33678", x"d6daa024", x"849ebb77", x"e92836bd"),
	(x"f8494430", x"cd130000", x"c3c80000", x"c6220000", x"a29461ae", x"45e0bb0c", x"1861ec49", x"a87a7517", x"e2cfa240", x"70de0000", x"5a8d0000", x"d0af0000", x"13bc0a7e", x"92df15dd", x"e28ab126", x"7b676bb7"),
	(x"17424640", x"f7ee0000", x"9e660000", x"af6b0000", x"399b5da8", x"01e50ef5", x"7e75e618", x"3a35281d", x"2ba4a270", x"97fb0000", x"75090000", x"f6e00000", x"1bd55187", x"ff23e4ea", x"b215d8a2", x"e50ec4df"),
	(x"25787800", x"93df0000", x"8d6b0000", x"110c0000", x"649c073b", x"98557743", x"0f57e2ed", x"d79dfeba", x"e7c8b400", x"65bf0000", x"dc600000", x"64dc0000", x"f31749e4", x"4380f45a", x"d6c5d8cc", x"ab657fca"),
	(x"ca737a70", x"a9220000", x"d0c50000", x"78450000", x"ff933b3d", x"dc50c2ba", x"6943e8bc", x"45d2a3b0", x"2ea3b430", x"829a0000", x"f3e40000", x"42930000", x"fb7e121d", x"2e7c056d", x"865ab148", x"350cd0a2"),
	(x"ec137830", x"74fa0000", x"a2ef0000", x"37430000", x"6cf55cc2", x"f5a98674", x"5fc88b69", x"49f451d2", x"c1a8b640", x"b8670000", x"ae4a0000", x"2bda0000", x"60712e1b", x"6a79b094", x"e04ebb19", x"a7438da8"),
	(x"03187a40", x"4e070000", x"ff410000", x"5e0a0000", x"f7fa60c4", x"b1ac338d", x"39dc8138", x"dbbb0cd8", x"08c3b670", x"5f420000", x"81ce0000", x"0d950000", x"681875e2", x"078541a3", x"b0d1d29d", x"392a22c0"),
	(x"dad61400", x"b8b10000", x"4f0c0000", x"574e0000", x"33a83a07", x"a50bfe67", x"628cfdb5", x"c7e6c5cb", x"a7bad400", x"36bb0000", x"78910000", x"34780000", x"8ed413f8", x"676c0dc3", x"fadcfe71", x"1ff06c8d"),
	(x"35dd1670", x"824c0000", x"12a20000", x"3e070000", x"a8a70601", x"e10e4b9e", x"0498f7e4", x"55a998c1", x"6ed1d430", x"d19e0000", x"57150000", x"12370000", x"86bd4801", x"0a90fcf4", x"aa4397f5", x"8199c3e5"),
	(x"13bd1430", x"5f940000", x"60880000", x"71010000", x"3bc161fe", x"c8f70f50", x"32139431", x"598f6aa3", x"81dad640", x"eb630000", x"0abb0000", x"7b7e0000", x"1db27407", x"4e95490d", x"cc579da4", x"13d69eef"),
	(x"fcb61640", x"65690000", x"3d260000", x"18480000", x"a0ce5df8", x"8cf2baa9", x"54079e60", x"cbc037a9", x"48b1d670", x"0c460000", x"253f0000", x"5d310000", x"15db2ffe", x"2369b83a", x"9cc8f420", x"8dbf3187"),
	(x"ce8c2800", x"01580000", x"2e2b0000", x"a62f0000", x"fdc9076b", x"1542c31f", x"25259a95", x"2668e10e", x"84ddc000", x"fe020000", x"8c560000", x"cf0d0000", x"fd19379d", x"9fcaa88a", x"f818f44e", x"c3d48a92"),
	(x"21872a70", x"3ba50000", x"73850000", x"cf660000", x"66c63b6d", x"514776e6", x"433190c4", x"b427bc04", x"4db6c030", x"19270000", x"a3d20000", x"e9420000", x"f5706c64", x"f23659bd", x"a8879dca", x"5dbd25fa"),
	(x"07e72830", x"e67d0000", x"01af0000", x"80600000", x"f5a05c92", x"78be3228", x"75baf311", x"b8014e66", x"a2bdc240", x"23da0000", x"fe7c0000", x"800b0000", x"6e7f5062", x"b633ec44", x"ce93979b", x"cff278f0"),
	(x"e8ec2a40", x"dc800000", x"5c010000", x"e9290000", x"6eaf6094", x"3cbb87d1", x"13aef940", x"2a4e136c", x"6bd6c270", x"c4ff0000", x"d1f80000", x"a6440000", x"66160b9b", x"dbcf1d73", x"9e0cfe1f", x"519bd798"),
	(x"f9b10000", x"70080000", x"bbcb0000", x"ac3b0000", x"40651e62", x"5dad5b2e", x"6048f78a", x"1bc223d4", x"9087fc00", x"47eb0000", x"ed710000", x"3e6c0000", x"33780af1", x"2f8395f2", x"bfb1936e", x"225aae57"),
	(x"16ba0270", x"4af50000", x"e6650000", x"c5720000", x"db6a2264", x"19a8eed7", x"065cfddb", x"898d7ede", x"59ecfc30", x"a0ce0000", x"c2f50000", x"18230000", x"3b115108", x"427f64c5", x"ef2efaea", x"bc33013f"),
	(x"30da0030", x"972d0000", x"944f0000", x"8a740000", x"480c459b", x"3051aa19", x"30d79e0e", x"85ab8cbc", x"b6e7fe40", x"9a330000", x"9f5b0000", x"716a0000", x"a01e6d0e", x"067ad13c", x"893af0bb", x"2e7c5c35"),
	(x"dfd10240", x"add00000", x"c9e10000", x"e33d0000", x"d303799d", x"74541fe0", x"56c3945f", x"17e4d1b6", x"7f8cfe70", x"7d160000", x"b0df0000", x"57250000", x"a87736f7", x"6b86200b", x"d9a5993f", x"b015f35d"),
	(x"edeb3c00", x"c9e10000", x"daec0000", x"5d5a0000", x"8e04230e", x"ede46656", x"27e190aa", x"fa4c0711", x"b3e0e800", x"8f520000", x"19b60000", x"c5190000", x"40b52e94", x"d72530bb", x"bd759951", x"fe7e4848"),
	(x"02e03e70", x"f31c0000", x"87420000", x"34130000", x"150b1f08", x"a9e1d3af", x"41f59afb", x"68035a1b", x"7a8be830", x"68770000", x"36320000", x"e3560000", x"48dc756d", x"bad9c18c", x"edeaf0d5", x"6017e720"),
	(x"24803c30", x"2ec40000", x"f5680000", x"7b150000", x"866d78f7", x"80189761", x"777ef92e", x"6425a879", x"9580ea40", x"528a0000", x"6b9c0000", x"8a1f0000", x"d3d3496b", x"fedc7475", x"8bfefa84", x"f258ba2a"),
	(x"cb8b3e40", x"14390000", x"a8c60000", x"125c0000", x"1d6244f1", x"c41d2298", x"116af37f", x"f66af573", x"5cebea70", x"b5af0000", x"44180000", x"ac500000", x"dbba1292", x"93208542", x"db619300", x"6c311542"),
	(x"8efe4800", x"525c0000", x"8ada0000", x"f68b0000", x"800a5d77", x"31ae3a86", x"093cbc28", x"92fdf249", x"3b01cc00", x"86680000", x"eac00000", x"d9eb0000", x"d7ee50bd", x"8678d837", x"b9dacdab", x"673aa2a4"),
	(x"61f54a70", x"68a10000", x"d7740000", x"9fc20000", x"1b056171", x"75ab8f7f", x"6f28b679", x"00b2af43", x"f26acc30", x"614d0000", x"c5440000", x"ffa40000", x"df870b44", x"eb842900", x"e945a42f", x"f9530dcc"),
	(x"47954830", x"b5790000", x"a55e0000", x"d0c40000", x"8863068e", x"5c52cbb1", x"59a3d5ac", x"0c945d21", x"1d61ce40", x"5bb00000", x"98ea0000", x"96ed0000", x"44883742", x"af819cf9", x"8f51ae7e", x"6b1c50c6"),
	(x"a89e4a40", x"8f840000", x"f8f00000", x"b98d0000", x"136c3a88", x"18577e48", x"3fb7dffd", x"9edb002b", x"d40ace70", x"bc950000", x"b76e0000", x"b0a20000", x"4ce16cbb", x"c27d6dce", x"dfcec7fa", x"f575ffae"),
	(x"9aa47400", x"ebb50000", x"ebfd0000", x"07ea0000", x"4e6b601b", x"81e707fe", x"4e95db08", x"7373d68c", x"1866d800", x"4ed10000", x"1e070000", x"229e0000", x"a42374d8", x"7ede7d7e", x"bb1ec794", x"bb1e44bb"),
	(x"75af7670", x"d1480000", x"b6530000", x"6ea30000", x"d5645c1d", x"c5e2b207", x"2881d159", x"e13c8b86", x"d10dd830", x"a9f40000", x"31830000", x"04d10000", x"ac4a2f21", x"13228c49", x"eb81ae10", x"2577ebd3"),
	(x"53cf7430", x"0c900000", x"c4790000", x"21a50000", x"46023be2", x"ec1bf6c9", x"1e0ab28c", x"ed1a79e4", x"3e06da40", x"93090000", x"6c2d0000", x"6d980000", x"37451327", x"572739b0", x"8d95a441", x"b738b6d9"),
	(x"bcc47640", x"366d0000", x"99d70000", x"48ec0000", x"dd0d07e4", x"a81e4330", x"781eb8dd", x"7f5524ee", x"f76dda70", x"742c0000", x"43a90000", x"4bd70000", x"3f2c48de", x"3adbc887", x"dd0acdc5", x"295119b1"),
	(x"ad995c00", x"9ae50000", x"7e1d0000", x"0dfe0000", x"f3c77912", x"c9089fcf", x"0bf8b617", x"4ed91456", x"0c3ce400", x"f7380000", x"7f200000", x"d3ff0000", x"6a4249b4", x"ce974006", x"fcb7a0b4", x"5a90607e"),
	(x"42925e70", x"a0180000", x"23b30000", x"64b70000", x"68c84514", x"8d0d2a36", x"6decbc46", x"dc96495c", x"c557e430", x"101d0000", x"50a40000", x"f5b00000", x"622b124d", x"a36bb131", x"ac28c930", x"c4f9cf16"),
	(x"64f25c30", x"7dc00000", x"51990000", x"2bb10000", x"fbae22eb", x"a4f46ef8", x"5b67df93", x"d0b0bb3e", x"2a5ce640", x"2ae00000", x"0d0a0000", x"9cf90000", x"f9242e4b", x"e76e04c8", x"ca3cc361", x"56b6921c"),
	(x"8bf95e40", x"473d0000", x"0c370000", x"42f80000", x"60a11eed", x"e0f1db01", x"3d73d5c2", x"42ffe634", x"e337e670", x"cdc50000", x"228e0000", x"bab60000", x"f14d75b2", x"8a92f5ff", x"9aa3aae5", x"c8df3d74"),
	(x"b9c36000", x"230c0000", x"1f3a0000", x"fc9f0000", x"3da6447e", x"7941a2b7", x"4c51d137", x"af573093", x"2f5bf000", x"3f810000", x"8be70000", x"288a0000", x"198f6dd1", x"3631e54f", x"fe73aa8b", x"86b48661"),
	(x"56c86270", x"19f10000", x"42940000", x"95d60000", x"a6a97878", x"3d44174e", x"2a45db66", x"3d186d99", x"e630f030", x"d8a40000", x"a4630000", x"0ec50000", x"11e63628", x"5bcd1478", x"aeecc30f", x"18dd2909"),
	(x"70a86030", x"c4290000", x"30be0000", x"dad00000", x"35cf1f87", x"14bd5380", x"1cceb8b3", x"313e9ffb", x"093bf240", x"e2590000", x"f9cd0000", x"678c0000", x"8ae90a2e", x"1fc8a181", x"c8f8c95e", x"8a927403"),
	(x"9fa36240", x"fed40000", x"6d100000", x"b3990000", x"aec02381", x"50b8e679", x"7adab2e2", x"a371c2f1", x"c050f270", x"057c0000", x"d6490000", x"41c30000", x"828051d7", x"723450b6", x"9867a0da", x"14fbdb6b"),
	(x"6f299000", x"6c850000", x"2f160000", x"782e0000", x"644c37cd", x"12dd1cd6", x"d26a8c36", x"32219526", x"29449c00", x"64e70000", x"f24b0000", x"c2f30000", x"0ede4e8f", x"56c23745", x"f3e04259", x"8d0d9ec4"),
	(x"80229270", x"56780000", x"72b80000", x"11670000", x"ff430bcb", x"56d8a92f", x"b47e8667", x"a06ec82c", x"e02f9c30", x"83c20000", x"ddcf0000", x"e4bc0000", x"06b71576", x"3b3ec672", x"a37f2bdd", x"136431ac"),
	(x"a6429030", x"8ba00000", x"00920000", x"5e610000", x"6c256c34", x"7f21ede1", x"82f5e5b2", x"ac483a4e", x"0f249e40", x"b93f0000", x"80610000", x"8df50000", x"9db82970", x"7f3b738b", x"c56b218c", x"812b6ca6"),
	(x"49499240", x"b15d0000", x"5d3c0000", x"37280000", x"f72a5032", x"3b245818", x"e4e1efe3", x"3e076744", x"c64f9e70", x"5e1a0000", x"afe50000", x"abba0000", x"95d17289", x"12c782bc", x"95f44808", x"1f42c3ce"),
	(x"7b73ac00", x"d56c0000", x"4e310000", x"894f0000", x"aa2d0aa1", x"a29421ae", x"95c3eb16", x"d3afb1e3", x"0a238800", x"ac5e0000", x"068c0000", x"39860000", x"7d136aea", x"ae64920c", x"f1244866", x"512978db"),
	(x"9478ae70", x"ef910000", x"139f0000", x"e0060000", x"312236a7", x"e6919457", x"f3d7e147", x"41e0ece9", x"c3488830", x"4b7b0000", x"29080000", x"1fc90000", x"757a3113", x"c398633b", x"a1bb21e2", x"cf40d7b3"),
	(x"b218ac30", x"32490000", x"61b50000", x"af000000", x"a2445158", x"cf68d099", x"c55c8292", x"4dc61e8b", x"2c438a40", x"71860000", x"74a60000", x"76800000", x"ee750d15", x"879dd6c2", x"c7af2bb3", x"5d0f8ab9"),
	(x"5d13ae40", x"08b40000", x"3c1b0000", x"c6490000", x"394b6d5e", x"8b6d6560", x"a34888c3", x"df894381", x"e5288a70", x"96a30000", x"5b220000", x"50cf0000", x"e61c56ec", x"ea6127f5", x"97304237", x"c36625d1"),
	(x"4c4e8400", x"a43c0000", x"dbd10000", x"835b0000", x"178113a8", x"ea7bb99f", x"d0ae8609", x"ee057339", x"1e79b400", x"15b70000", x"67ab0000", x"c8e70000", x"b3725786", x"1e2daf74", x"b68d2f46", x"b0a75c1e"),
	(x"a3458670", x"9ec10000", x"867f0000", x"ea120000", x"8c8e2fae", x"ae7e0c66", x"b6ba8c58", x"7c4a2e33", x"d712b430", x"f2920000", x"482f0000", x"eea80000", x"bb1b0c7f", x"73d15e43", x"e61246c2", x"2ecef376"),
	(x"85258430", x"43190000", x"f4550000", x"a5140000", x"1fe84851", x"878748a8", x"8031ef8d", x"706cdc51", x"3819b640", x"c86f0000", x"15810000", x"87e10000", x"20143079", x"37d4ebba", x"80064c93", x"bc81ae7c"),
	(x"6a2e8640", x"79e40000", x"a9fb0000", x"cc5d0000", x"84e77457", x"c382fd51", x"e625e5dc", x"e223815b", x"f172b670", x"2f4a0000", x"3a050000", x"a1ae0000", x"287d6b80", x"5a281a8d", x"d0992517", x"22e80114"),
	(x"5814b800", x"1dd50000", x"baf60000", x"723a0000", x"d9e02ec4", x"5a3284e7", x"9707e129", x"0f8b57fc", x"3d1ea000", x"dd0e0000", x"936c0000", x"33920000", x"c0bf73e3", x"e68b0a3d", x"b4492579", x"6c83ba01"),
	(x"b71fba70", x"27280000", x"e7580000", x"1b730000", x"42ef12c2", x"1e37311e", x"f113eb78", x"9dc40af6", x"f475a030", x"3a2b0000", x"bce80000", x"15dd0000", x"c8d6281a", x"8b77fb0a", x"e4d64cfd", x"f2ea1569"),
	(x"917fb830", x"faf00000", x"95720000", x"54750000", x"d189753d", x"37ce75d0", x"c79888ad", x"91e2f894", x"1b7ea240", x"00d60000", x"e1460000", x"7c940000", x"53d9141c", x"cf724ef3", x"82c246ac", x"60a54863"),
	(x"7e74ba40", x"c00d0000", x"c8dc0000", x"3d3c0000", x"4a86493b", x"73cbc029", x"a18c82fc", x"03ada59e", x"d215a270", x"e7f30000", x"cec20000", x"5adb0000", x"5bb04fe5", x"a28ebfc4", x"d25d2f28", x"fecce70b"),
	(x"3b01cc00", x"86680000", x"eac00000", x"d9eb0000", x"d7ee50bd", x"8678d837", x"b9dacdab", x"673aa2a4", x"b5ff8400", x"d4340000", x"601a0000", x"2f600000", x"57e40dca", x"b7d6e2b1", x"b0e67183", x"f5c750ed"),
	(x"d40ace70", x"bc950000", x"b76e0000", x"b0a20000", x"4ce16cbb", x"c27d6dce", x"dfcec7fa", x"f575ffae", x"7c948430", x"33110000", x"4f9e0000", x"092f0000", x"5f8d5633", x"da2a1386", x"e0791807", x"6baeff85"),
	(x"f26acc30", x"614d0000", x"c5440000", x"ffa40000", x"df870b44", x"eb842900", x"e945a42f", x"f9530dcc", x"939f8640", x"09ec0000", x"12300000", x"60660000", x"c4826a35", x"9e2fa67f", x"866d1256", x"f9e1a28f"),
	(x"1d61ce40", x"5bb00000", x"98ea0000", x"96ed0000", x"44883742", x"af819cf9", x"8f51ae7e", x"6b1c50c6", x"5af48670", x"eec90000", x"3db40000", x"46290000", x"cceb31cc", x"f3d35748", x"d6f27bd2", x"67880de7"),
	(x"2f5bf000", x"3f810000", x"8be70000", x"288a0000", x"198f6dd1", x"3631e54f", x"fe73aa8b", x"86b48661", x"96989000", x"1c8d0000", x"94dd0000", x"d4150000", x"242929af", x"4f7047f8", x"b2227bbc", x"29e3b6f2"),
	(x"c050f270", x"057c0000", x"d6490000", x"41c30000", x"828051d7", x"723450b6", x"9867a0da", x"14fbdb6b", x"5ff39030", x"fba80000", x"bb590000", x"f25a0000", x"2c407256", x"228cb6cf", x"e2bd1238", x"b78a199a"),
	(x"e630f030", x"d8a40000", x"a4630000", x"0ec50000", x"11e63628", x"5bcd1478", x"aeecc30f", x"18dd2909", x"b0f89240", x"c1550000", x"e6f70000", x"9b130000", x"b74f4e50", x"66890336", x"84a91869", x"25c54490"),
	(x"093bf240", x"e2590000", x"f9cd0000", x"678c0000", x"8ae90a2e", x"1fc8a181", x"c8f8c95e", x"8a927403", x"79939270", x"26700000", x"c9730000", x"bd5c0000", x"bf2615a9", x"0b75f201", x"d43671ed", x"bbacebf8"),
	(x"1866d800", x"4ed10000", x"1e070000", x"229e0000", x"a42374d8", x"7ede7d7e", x"bb1ec794", x"bb1e44bb", x"82c2ac00", x"a5640000", x"f5fa0000", x"25740000", x"ea4814c3", x"ff397a80", x"f58b1c9c", x"c86d9237"),
	(x"f76dda70", x"742c0000", x"43a90000", x"4bd70000", x"3f2c48de", x"3adbc887", x"dd0acdc5", x"295119b1", x"4ba9ac30", x"42410000", x"da7e0000", x"033b0000", x"e2214f3a", x"92c58bb7", x"a5147518", x"56043d5f"),
	(x"d10dd830", x"a9f40000", x"31830000", x"04d10000", x"ac4a2f21", x"13228c49", x"eb81ae10", x"2577ebd3", x"a4a2ae40", x"78bc0000", x"87d00000", x"6a720000", x"792e733c", x"d6c03e4e", x"c3007f49", x"c44b6055"),
	(x"3e06da40", x"93090000", x"6c2d0000", x"6d980000", x"37451327", x"572739b0", x"8d95a441", x"b738b6d9", x"6dc9ae70", x"9f990000", x"a8540000", x"4c3d0000", x"714728c5", x"bb3ccf79", x"939f16cd", x"5a22cf3d"),
	(x"0c3ce400", x"f7380000", x"7f200000", x"d3ff0000", x"6a4249b4", x"ce974006", x"fcb7a0b4", x"5a90607e", x"a1a5b800", x"6ddd0000", x"013d0000", x"de010000", x"998530a6", x"079fdfc9", x"f74f16a3", x"14497428"),
	(x"e337e670", x"cdc50000", x"228e0000", x"bab60000", x"f14d75b2", x"8a92f5ff", x"9aa3aae5", x"c8df3d74", x"68ceb830", x"8af80000", x"2eb90000", x"f84e0000", x"91ec6b5f", x"6a632efe", x"a7d07f27", x"8a20db40"),
	(x"c557e430", x"101d0000", x"50a40000", x"f5b00000", x"622b124d", x"a36bb131", x"ac28c930", x"c4f9cf16", x"87c5ba40", x"b0050000", x"73170000", x"91070000", x"0ae35759", x"2e669b07", x"c1c47576", x"186f864a"),
	(x"2a5ce640", x"2ae00000", x"0d0a0000", x"9cf90000", x"f9242e4b", x"e76e04c8", x"ca3cc361", x"56b6921c", x"4eaeba70", x"57200000", x"5c930000", x"b7480000", x"028a0ca0", x"439a6a30", x"915b1cf2", x"86062922"),
	(x"f3928800", x"dc560000", x"bd470000", x"95bd0000", x"3d767488", x"f3c9c922", x"916cbfec", x"4aeb5b0f", x"e1d7d800", x"3ed90000", x"a5cc0000", x"8ea50000", x"e4466aba", x"23732650", x"db56301e", x"a0dc676f"),
	(x"1c998a70", x"e6ab0000", x"e0e90000", x"fcf40000", x"a679488e", x"b7cc7cdb", x"f778b5bd", x"d8a40605", x"28bcd830", x"d9fc0000", x"8a480000", x"a8ea0000", x"ec2f3143", x"4e8fd767", x"8bc9599a", x"3eb5c807"),
	(x"3af98830", x"3b730000", x"92c30000", x"b3f20000", x"351f2f71", x"9e353815", x"c1f3d668", x"d482f467", x"c7b7da40", x"e3010000", x"d7e60000", x"c1a30000", x"77200d45", x"0a8a629e", x"eddd53cb", x"acfa950d"),
	(x"d5f28a40", x"018e0000", x"cf6d0000", x"dabb0000", x"ae101377", x"da308dec", x"a7e7dc39", x"46cda96d", x"0edcda70", x"04240000", x"f8620000", x"e7ec0000", x"7f4956bc", x"677693a9", x"bd423a4f", x"32933a65"),
	(x"e7c8b400", x"65bf0000", x"dc600000", x"64dc0000", x"f31749e4", x"4380f45a", x"d6c5d8cc", x"ab657fca", x"c2b0cc00", x"f6600000", x"510b0000", x"75d00000", x"978b4edf", x"dbd58319", x"d9923a21", x"7cf88170"),
	(x"08c3b670", x"5f420000", x"81ce0000", x"0d950000", x"681875e2", x"078541a3", x"b0d1d29d", x"392a22c0", x"0bdbcc30", x"11450000", x"7e8f0000", x"539f0000", x"9fe21526", x"b629722e", x"890d53a5", x"e2912e18"),
	(x"2ea3b430", x"829a0000", x"f3e40000", x"42930000", x"fb7e121d", x"2e7c056d", x"865ab148", x"350cd0a2", x"e4d0ce40", x"2bb80000", x"23210000", x"3ad60000", x"04ed2920", x"f22cc7d7", x"ef1959f4", x"70de7312"),
	(x"c1a8b640", x"b8670000", x"ae4a0000", x"2bda0000", x"60712e1b", x"6a79b094", x"e04ebb19", x"a7438da8", x"2dbbce70", x"cc9d0000", x"0ca50000", x"1c990000", x"0c8472d9", x"9fd036e0", x"bf863070", x"eeb7dc7a"),
	(x"d0f59c00", x"14ef0000", x"49800000", x"6ec80000", x"4ebb50ed", x"0b6f6c6b", x"93a8b5d3", x"96cfbd10", x"d6eaf000", x"4f890000", x"302c0000", x"84b10000", x"59ea73b3", x"6b9cbe61", x"9e3b5d01", x"9d76a5b5"),
	(x"3ffe9e70", x"2e120000", x"142e0000", x"07810000", x"d5b46ceb", x"4f6ad992", x"f5bcbf82", x"0480e01a", x"1f81f030", x"a8ac0000", x"1fa80000", x"a2fe0000", x"5183284a", x"06604f56", x"cea43485", x"031f0add"),
	(x"199e9c30", x"f3ca0000", x"66040000", x"48870000", x"46d20b14", x"66939d5c", x"c337dc57", x"08a61278", x"f08af240", x"92510000", x"42060000", x"cbb70000", x"ca8c144c", x"4265faaf", x"a8b03ed4", x"915057d7"),
	(x"f6959e40", x"c9370000", x"3baa0000", x"21ce0000", x"dddd3712", x"229628a5", x"a523d606", x"9ae94f72", x"39e1f270", x"75740000", x"6d820000", x"edf80000", x"c2e54fb5", x"2f990b98", x"f82f5750", x"0f39f8bf"),
	(x"c4afa000", x"ad060000", x"28a70000", x"9fa90000", x"80da6d81", x"bb265113", x"d401d2f3", x"774199d5", x"f58de400", x"87300000", x"c4eb0000", x"7fc40000", x"2a2757d6", x"933a1b28", x"9cff573e", x"415243aa"),
	(x"2ba4a270", x"97fb0000", x"75090000", x"f6e00000", x"1bd55187", x"ff23e4ea", x"b215d8a2", x"e50ec4df", x"3ce6e430", x"60150000", x"eb6f0000", x"598b0000", x"224e0c2f", x"fec6ea1f", x"cc603eba", x"df3becc2"),
	(x"0dc4a030", x"4a230000", x"07230000", x"b9e60000", x"88b33678", x"d6daa024", x"849ebb77", x"e92836bd", x"d3ede640", x"5ae80000", x"b6c10000", x"30c20000", x"b9413029", x"bac35fe6", x"aa7434eb", x"4d74b1c8"),
	(x"e2cfa240", x"70de0000", x"5a8d0000", x"d0af0000", x"13bc0a7e", x"92df15dd", x"e28ab126", x"7b676bb7", x"1a86e670", x"bdcd0000", x"99450000", x"168d0000", x"b1286bd0", x"d73faed1", x"faeb5d6f", x"d31d1ea0"),
	(x"a7bad400", x"36bb0000", x"78910000", x"34780000", x"8ed413f8", x"676c0dc3", x"fadcfe71", x"1ff06c8d", x"7d6cc000", x"8e0a0000", x"379d0000", x"63360000", x"bd7c29ff", x"c267f3a4", x"985003c4", x"d816a946"),
	(x"48b1d670", x"0c460000", x"253f0000", x"5d310000", x"15db2ffe", x"2369b83a", x"9cc8f420", x"8dbf3187", x"b407c030", x"692f0000", x"18190000", x"45790000", x"b5157206", x"af9b0293", x"c8cf6a40", x"467f062e"),
	(x"6ed1d430", x"d19e0000", x"57150000", x"12370000", x"86bd4801", x"0a90fcf4", x"aa4397f5", x"8199c3e5", x"5b0cc240", x"53d20000", x"45b70000", x"2c300000", x"2e1a4e00", x"eb9eb76a", x"aedb6011", x"d4305b24"),
	(x"81dad640", x"eb630000", x"0abb0000", x"7b7e0000", x"1db27407", x"4e95490d", x"cc579da4", x"13d69eef", x"9267c270", x"b4f70000", x"6a330000", x"0a7f0000", x"267315f9", x"8662465d", x"fe440995", x"4a59f44c"),
	(x"b3e0e800", x"8f520000", x"19b60000", x"c5190000", x"40b52e94", x"d72530bb", x"bd759951", x"fe7e4848", x"5e0bd400", x"46b30000", x"c35a0000", x"98430000", x"ceb10d9a", x"3ac156ed", x"9a9409fb", x"04324f59"),
	(x"5cebea70", x"b5af0000", x"44180000", x"ac500000", x"dbba1292", x"93208542", x"db619300", x"6c311542", x"9760d430", x"a1960000", x"ecde0000", x"be0c0000", x"c6d85663", x"573da7da", x"ca0b607f", x"9a5be031"),
	(x"7a8be830", x"68770000", x"36320000", x"e3560000", x"48dc756d", x"bad9c18c", x"edeaf0d5", x"6017e720", x"786bd640", x"9b6b0000", x"b1700000", x"d7450000", x"5dd76a65", x"13381223", x"ac1f6a2e", x"0814bd3b"),
	(x"9580ea40", x"528a0000", x"6b9c0000", x"8a1f0000", x"d3d3496b", x"fedc7475", x"8bfefa84", x"f258ba2a", x"b100d670", x"7c4e0000", x"9ef40000", x"f10a0000", x"55be319c", x"7ec4e314", x"fc8003aa", x"967d1253"),
	(x"84ddc000", x"fe020000", x"8c560000", x"cf0d0000", x"fd19379d", x"9fcaa88a", x"f818f44e", x"c3d48a92", x"4a51e800", x"ff5a0000", x"a27d0000", x"69220000", x"00d030f6", x"8a886b95", x"dd3d6edb", x"e5bc6b9c"),
	(x"6bd6c270", x"c4ff0000", x"d1f80000", x"a6440000", x"66160b9b", x"dbcf1d73", x"9e0cfe1f", x"519bd798", x"833ae830", x"187f0000", x"8df90000", x"4f6d0000", x"08b96b0f", x"e7749aa2", x"8da2075f", x"7bd5c4f4"),
	(x"4db6c030", x"19270000", x"a3d20000", x"e9420000", x"f5706c64", x"f23659bd", x"a8879dca", x"5dbd25fa", x"6c31ea40", x"22820000", x"d0570000", x"26240000", x"93b65709", x"a3712f5b", x"ebb60d0e", x"e99a99fe"),
	(x"a2bdc240", x"23da0000", x"fe7c0000", x"800b0000", x"6e7f5062", x"b633ec44", x"ce93979b", x"cff278f0", x"a55aea70", x"c5a70000", x"ffd30000", x"006b0000", x"9bdf0cf0", x"ce8dde6c", x"bb29648a", x"77f33696"),
	(x"9087fc00", x"47eb0000", x"ed710000", x"3e6c0000", x"33780af1", x"2f8395f2", x"bfb1936e", x"225aae57", x"6936fc00", x"37e30000", x"56ba0000", x"92570000", x"731d1493", x"722ecedc", x"dff964e4", x"39988d83"),
	(x"7f8cfe70", x"7d160000", x"b0df0000", x"57250000", x"a87736f7", x"6b86200b", x"d9a5993f", x"b015f35d", x"a05dfc30", x"d0c60000", x"793e0000", x"b4180000", x"7b744f6a", x"1fd23feb", x"8f660d60", x"a7f122eb"),
	(x"59ecfc30", x"a0ce0000", x"c2f50000", x"18230000", x"3b115108", x"427f64c5", x"ef2efaea", x"bc33013f", x"4f56fe40", x"ea3b0000", x"24900000", x"dd510000", x"e07b736c", x"5bd78a12", x"e9720731", x"35be7fe1"),
	(x"b6e7fe40", x"9a330000", x"9f5b0000", x"716a0000", x"a01e6d0e", x"067ad13c", x"893af0bb", x"2e7c5c35", x"863dfe70", x"0d1e0000", x"0b140000", x"fb1e0000", x"e8122895", x"362b7b25", x"b9ed6eb5", x"abd7d089")
    ),(
	(x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000"),
	(x"f6800005", x"3443c000", x"24070000", x"8f3d0000", x"21373bfb", x"0ab8d5ae", x"cdc58b19", x"d795ba31", x"a67f0001", x"71378000", x"19fc0000", x"96db0000", x"3a8b6dfd", x"ebcaaef3", x"2c6d478f", x"ac8e6c88"),
	(x"a67f0001", x"71378000", x"19fc0000", x"96db0000", x"3a8b6dfd", x"ebcaaef3", x"2c6d478f", x"ac8e6c88", x"50ff0004", x"45744000", x"3dfb0000", x"19e60000", x"1bbc5606", x"e1727b5d", x"e1a8cc96", x"7b1bd6b9"),
	(x"50ff0004", x"45744000", x"3dfb0000", x"19e60000", x"1bbc5606", x"e1727b5d", x"e1a8cc96", x"7b1bd6b9", x"f6800005", x"3443c000", x"24070000", x"8f3d0000", x"21373bfb", x"0ab8d5ae", x"cdc58b19", x"d795ba31"),
	(x"f7750009", x"cf3cc000", x"c3d60000", x"04920000", x"029519a9", x"f8e836ba", x"7a87f14e", x"9e16981a", x"d46a0000", x"8dc8c000", x"a5af0000", x"4a290000", x"fc4e427a", x"c9b4866c", x"98369604", x"f746c320"),
	(x"01f5000c", x"fb7f0000", x"e7d10000", x"8baf0000", x"23a22252", x"f250e314", x"b7427a57", x"4983222b", x"72150001", x"fcff4000", x"bc530000", x"dcf20000", x"c6c52f87", x"227e289f", x"b45bd18b", x"5bc8afa8"),
	(x"510a0008", x"be0b4000", x"da2a0000", x"92490000", x"381e7454", x"13229849", x"56eab6c1", x"3298f492", x"84950004", x"c8bc8000", x"98540000", x"53cf0000", x"e7f2147c", x"28c6fd31", x"799e5a92", x"8c5d1599"),
	(x"a78a000d", x"8a488000", x"fe2d0000", x"1d740000", x"19294faf", x"199a4de7", x"9b2f3dd8", x"e50d4ea3", x"22ea0005", x"b98b0000", x"81a80000", x"c5140000", x"dd797981", x"c30c53c2", x"55f31d1d", x"20d37911"),
	(x"d46a0000", x"8dc8c000", x"a5af0000", x"4a290000", x"fc4e427a", x"c9b4866c", x"98369604", x"f746c320", x"231f0009", x"42f40000", x"66790000", x"4ebb0000", x"fedb5bd3", x"315cb0d6", x"e2b1674a", x"69505b3a"),
	(x"22ea0005", x"b98b0000", x"81a80000", x"c5140000", x"dd797981", x"c30c53c2", x"55f31d1d", x"20d37911", x"85600008", x"33c38000", x"7f850000", x"d8600000", x"c450362e", x"da961e25", x"cedc20c5", x"c5de37b2"),
	(x"72150001", x"fcff4000", x"bc530000", x"dcf20000", x"c6c52f87", x"227e289f", x"b45bd18b", x"5bc8afa8", x"73e0000d", x"07804000", x"5b820000", x"575d0000", x"e5670dd5", x"d02ecb8b", x"0319abdc", x"124b8d83"),
	(x"84950004", x"c8bc8000", x"98540000", x"53cf0000", x"e7f2147c", x"28c6fd31", x"799e5a92", x"8c5d1599", x"d59f000c", x"76b7c000", x"427e0000", x"c1860000", x"dfec6028", x"3be46578", x"2f74ec53", x"bec5e10b"),
	(x"231f0009", x"42f40000", x"66790000", x"4ebb0000", x"fedb5bd3", x"315cb0d6", x"e2b1674a", x"69505b3a", x"f7750009", x"cf3cc000", x"c3d60000", x"04920000", x"029519a9", x"f8e836ba", x"7a87f14e", x"9e16981a"),
	(x"d59f000c", x"76b7c000", x"427e0000", x"c1860000", x"dfec6028", x"3be46578", x"2f74ec53", x"bec5e10b", x"510a0008", x"be0b4000", x"da2a0000", x"92490000", x"381e7454", x"13229849", x"56eab6c1", x"3298f492"),
	(x"85600008", x"33c38000", x"7f850000", x"d8600000", x"c450362e", x"da961e25", x"cedc20c5", x"c5de37b2", x"a78a000d", x"8a488000", x"fe2d0000", x"1d740000", x"19294faf", x"199a4de7", x"9b2f3dd8", x"e50d4ea3"),
	(x"73e0000d", x"07804000", x"5b820000", x"575d0000", x"e5670dd5", x"d02ecb8b", x"0319abdc", x"124b8d83", x"01f5000c", x"fb7f0000", x"e7d10000", x"8baf0000", x"23a22252", x"f250e314", x"b7427a57", x"4983222b"),
	(x"774400f0", x"f15a0000", x"f5b20000", x"34140000", x"89377e8c", x"5a8bec25", x"0bc3cd1e", x"cf3775cb", x"f46c0050", x"96180000", x"14a50000", x"031f0000", x"42947eb8", x"66bf7e19", x"9ca470d2", x"8a341574"),
	(x"81c400f5", x"c519c000", x"d1b50000", x"bb290000", x"a8004577", x"5033398b", x"c6064607", x"18a2cffa", x"52130051", x"e72f8000", x"0d590000", x"95c40000", x"781f1345", x"8d75d0ea", x"b0c9375d", x"26ba79fc"),
	(x"d13b00f1", x"806d8000", x"ec4e0000", x"a2cf0000", x"b3bc1371", x"b14142d6", x"27ae8a91", x"63b91943", x"a4930054", x"d36c4000", x"295e0000", x"1af90000", x"592828be", x"87cd0544", x"7d0cbc44", x"f12fc3cd"),
	(x"27bb00f4", x"b42e4000", x"c8490000", x"2df20000", x"928b288a", x"bbf99778", x"ea6b0188", x"b42ca372", x"02ec0055", x"a25bc000", x"30a20000", x"8c220000", x"63a34543", x"6c07abb7", x"5161fbcb", x"5da1af45"),
	(x"803100f9", x"3e66c000", x"36640000", x"30860000", x"8ba26725", x"a263da9f", x"71443c50", x"5121edd1", x"20060050", x"1bd0c000", x"b10a0000", x"49360000", x"beda3cc2", x"af0bf875", x"0492e6d6", x"7d72d654"),
	(x"76b100fc", x"0a250000", x"12630000", x"bfbb0000", x"aa955cde", x"a8db0f31", x"bc81b749", x"86b457e0", x"86790051", x"6ae74000", x"a8f60000", x"dfed0000", x"8451513f", x"44c15686", x"28ffa159", x"d1fcbadc"),
	(x"264e00f8", x"4f514000", x"2f980000", x"a65d0000", x"b1290ad8", x"49a9746c", x"5d297bdf", x"fdaf8159", x"70f90054", x"5ea48000", x"8cf10000", x"50d00000", x"a5666ac4", x"4e798328", x"e53a2a40", x"066900ed"),
	(x"d0ce00fd", x"7b128000", x"0b9f0000", x"29600000", x"901e3123", x"4311a1c2", x"90ecf0c6", x"2a3a3b68", x"d6860055", x"2f930000", x"950d0000", x"c60b0000", x"9fed0739", x"a5b32ddb", x"c9576dcf", x"aae76c65"),
	(x"a32e00f0", x"7c92c000", x"501d0000", x"7e3d0000", x"75793cf6", x"933f6a49", x"93f55b1a", x"3871b6eb", x"d7730059", x"d4ec0000", x"72dc0000", x"4da40000", x"bc4f256b", x"57e3cecf", x"7e151798", x"e3644e4e"),
	(x"55ae00f5", x"48d10000", x"741a0000", x"f1000000", x"544e070d", x"9987bfe7", x"5e30d003", x"efe40cda", x"710c0058", x"a5db8000", x"6b200000", x"db7f0000", x"86c44896", x"bc29603c", x"52785017", x"4fea22c6"),
	(x"055100f1", x"0da54000", x"49e10000", x"e8e60000", x"4ff2510b", x"78f5c4ba", x"bf981c95", x"94ffda63", x"878c005d", x"91984000", x"4f270000", x"54420000", x"a7f3736d", x"b691b592", x"9fbddb0e", x"987f98f7"),
	(x"f3d100f4", x"39e68000", x"6de60000", x"67db0000", x"6ec56af0", x"724d1114", x"725d978c", x"436a6052", x"21f3005c", x"e0afc000", x"56db0000", x"c2990000", x"9d781e90", x"5d5b1b61", x"b3d09c81", x"34f1f47f"),
	(x"545b00f9", x"b3ae0000", x"93cb0000", x"7aaf0000", x"77ec255f", x"6bd75cf3", x"e972aa54", x"a6672ef1", x"03190059", x"5924c000", x"d7730000", x"078d0000", x"40016711", x"9e5748a3", x"e623819c", x"14228d6e"),
	(x"a2db00fc", x"87edc000", x"b7cc0000", x"f5920000", x"56db1ea4", x"616f895d", x"24b7214d", x"71f294c0", x"a5660058", x"28134000", x"ce8f0000", x"91560000", x"7a8a0aec", x"759de650", x"ca4ec613", x"b8ace1e6"),
	(x"f22400f8", x"c2998000", x"8a370000", x"ec740000", x"4d6748a2", x"801df200", x"c51feddb", x"0ae94279", x"53e6005d", x"1c508000", x"ea880000", x"1e6b0000", x"5bbd3117", x"7f2533fe", x"078b4d0a", x"6f395bd7"),
	(x"04a400fd", x"f6da4000", x"ae300000", x"63490000", x"6c507359", x"8aa527ae", x"08da66c2", x"dd7cf848", x"f599005c", x"6d670000", x"f3740000", x"88b00000", x"61365cea", x"94ef9d0d", x"2be60a85", x"c3b7375f"),
	(x"f46c0050", x"96180000", x"14a50000", x"031f0000", x"42947eb8", x"66bf7e19", x"9ca470d2", x"8a341574", x"832800a0", x"67420000", x"e1170000", x"370b0000", x"cba30034", x"3c34923c", x"9767bdcc", x"450360bf"),
	(x"02ec0055", x"a25bc000", x"30a20000", x"8c220000", x"63a34543", x"6c07abb7", x"5161fbcb", x"5da1af45", x"255700a1", x"16758000", x"f8eb0000", x"a1d00000", x"f1286dc9", x"d7fe3ccf", x"bb0afa43", x"e98d0c37"),
	(x"52130051", x"e72f8000", x"0d590000", x"95c40000", x"781f1345", x"8d75d0ea", x"b0c9375d", x"26ba79fc", x"d3d700a4", x"22364000", x"dcec0000", x"2eed0000", x"d01f5632", x"dd46e961", x"76cf715a", x"3e18b606"),
	(x"a4930054", x"d36c4000", x"295e0000", x"1af90000", x"592828be", x"87cd0544", x"7d0cbc44", x"f12fc3cd", x"75a800a5", x"5301c000", x"c5100000", x"b8360000", x"ea943bcf", x"368c4792", x"5aa236d5", x"9296da8e"),
	(x"03190059", x"5924c000", x"d7730000", x"078d0000", x"40016711", x"9e5748a3", x"e623819c", x"14228d6e", x"574200a0", x"ea8ac000", x"44b80000", x"7d220000", x"37ed424e", x"f5801450", x"0f512bc8", x"b245a39f"),
	(x"f599005c", x"6d670000", x"f3740000", x"88b00000", x"61365cea", x"94ef9d0d", x"2be60a85", x"c3b7375f", x"f13d00a1", x"9bbd4000", x"5d440000", x"ebf90000", x"0d662fb3", x"1e4abaa3", x"233c6c47", x"1ecbcf17"),
	(x"a5660058", x"28134000", x"ce8f0000", x"91560000", x"7a8a0aec", x"759de650", x"ca4ec613", x"b8ace1e6", x"07bd00a4", x"affe8000", x"79430000", x"64c40000", x"2c511448", x"14f26f0d", x"eef9e75e", x"c95e7526"),
	(x"53e6005d", x"1c508000", x"ea880000", x"1e6b0000", x"5bbd3117", x"7f2533fe", x"078b4d0a", x"6f395bd7", x"a1c200a5", x"dec90000", x"60bf0000", x"f21f0000", x"16da79b5", x"ff38c1fe", x"c294a0d1", x"65d019ae"),
	(x"20060050", x"1bd0c000", x"b10a0000", x"49360000", x"beda3cc2", x"af0bf875", x"0492e6d6", x"7d72d654", x"a03700a9", x"25b60000", x"876e0000", x"79b00000", x"35785be7", x"0d6822ea", x"75d6da86", x"2c533b85"),
	(x"d6860055", x"2f930000", x"950d0000", x"c60b0000", x"9fed0739", x"a5b32ddb", x"c9576dcf", x"aae76c65", x"064800a8", x"54818000", x"9e920000", x"ef6b0000", x"0ff3361a", x"e6a28c19", x"59bb9d09", x"80dd570d"),
	(x"86790051", x"6ae74000", x"a8f60000", x"dfed0000", x"8451513f", x"44c15686", x"28ffa159", x"d1fcbadc", x"f0c800ad", x"60c24000", x"ba950000", x"60560000", x"2ec40de1", x"ec1a59b7", x"947e1610", x"5748ed3c"),
	(x"70f90054", x"5ea48000", x"8cf10000", x"50d00000", x"a5666ac4", x"4e798328", x"e53a2a40", x"066900ed", x"56b700ac", x"11f5c000", x"a3690000", x"f68d0000", x"144f601c", x"07d0f744", x"b813519f", x"fbc681b4"),
	(x"d7730059", x"d4ec0000", x"72dc0000", x"4da40000", x"bc4f256b", x"57e3cecf", x"7e151798", x"e3644e4e", x"745d00a9", x"a87ec000", x"22c10000", x"33990000", x"c936199d", x"c4dca486", x"ede04c82", x"db15f8a5"),
	(x"21f3005c", x"e0afc000", x"56db0000", x"c2990000", x"9d781e90", x"5d5b1b61", x"b3d09c81", x"34f1f47f", x"d22200a8", x"d9494000", x"3b3d0000", x"a5420000", x"f3bd7460", x"2f160a75", x"c18d0b0d", x"779b942d"),
	(x"710c0058", x"a5db8000", x"6b200000", x"db7f0000", x"86c44896", x"bc29603c", x"52785017", x"4fea22c6", x"24a200ad", x"ed0a8000", x"1f3a0000", x"2a7f0000", x"d28a4f9b", x"25aedfdb", x"0c488014", x"a00e2e1c"),
	(x"878c005d", x"91984000", x"4f270000", x"54420000", x"a7f3736d", x"b691b592", x"9fbddb0e", x"987f98f7", x"82dd00ac", x"9c3d0000", x"06c60000", x"bca40000", x"e8012266", x"ce647128", x"2025c79b", x"0c804294"),
	(x"832800a0", x"67420000", x"e1170000", x"370b0000", x"cba30034", x"3c34923c", x"9767bdcc", x"450360bf", x"774400f0", x"f15a0000", x"f5b20000", x"34140000", x"89377e8c", x"5a8bec25", x"0bc3cd1e", x"cf3775cb"),
	(x"75a800a5", x"5301c000", x"c5100000", x"b8360000", x"ea943bcf", x"368c4792", x"5aa236d5", x"9296da8e", x"d13b00f1", x"806d8000", x"ec4e0000", x"a2cf0000", x"b3bc1371", x"b14142d6", x"27ae8a91", x"63b91943"),
	(x"255700a1", x"16758000", x"f8eb0000", x"a1d00000", x"f1286dc9", x"d7fe3ccf", x"bb0afa43", x"e98d0c37", x"27bb00f4", x"b42e4000", x"c8490000", x"2df20000", x"928b288a", x"bbf99778", x"ea6b0188", x"b42ca372"),
	(x"d3d700a4", x"22364000", x"dcec0000", x"2eed0000", x"d01f5632", x"dd46e961", x"76cf715a", x"3e18b606", x"81c400f5", x"c519c000", x"d1b50000", x"bb290000", x"a8004577", x"5033398b", x"c6064607", x"18a2cffa"),
	(x"745d00a9", x"a87ec000", x"22c10000", x"33990000", x"c936199d", x"c4dca486", x"ede04c82", x"db15f8a5", x"a32e00f0", x"7c92c000", x"501d0000", x"7e3d0000", x"75793cf6", x"933f6a49", x"93f55b1a", x"3871b6eb"),
	(x"82dd00ac", x"9c3d0000", x"06c60000", x"bca40000", x"e8012266", x"ce647128", x"2025c79b", x"0c804294", x"055100f1", x"0da54000", x"49e10000", x"e8e60000", x"4ff2510b", x"78f5c4ba", x"bf981c95", x"94ffda63"),
	(x"d22200a8", x"d9494000", x"3b3d0000", x"a5420000", x"f3bd7460", x"2f160a75", x"c18d0b0d", x"779b942d", x"f3d100f4", x"39e68000", x"6de60000", x"67db0000", x"6ec56af0", x"724d1114", x"725d978c", x"436a6052"),
	(x"24a200ad", x"ed0a8000", x"1f3a0000", x"2a7f0000", x"d28a4f9b", x"25aedfdb", x"0c488014", x"a00e2e1c", x"55ae00f5", x"48d10000", x"741a0000", x"f1000000", x"544e070d", x"9987bfe7", x"5e30d003", x"efe40cda"),
	(x"574200a0", x"ea8ac000", x"44b80000", x"7d220000", x"37ed424e", x"f5801450", x"0f512bc8", x"b245a39f", x"545b00f9", x"b3ae0000", x"93cb0000", x"7aaf0000", x"77ec255f", x"6bd75cf3", x"e972aa54", x"a6672ef1"),
	(x"a1c200a5", x"dec90000", x"60bf0000", x"f21f0000", x"16da79b5", x"ff38c1fe", x"c294a0d1", x"65d019ae", x"f22400f8", x"c2998000", x"8a370000", x"ec740000", x"4d6748a2", x"801df200", x"c51feddb", x"0ae94279"),
	(x"f13d00a1", x"9bbd4000", x"5d440000", x"ebf90000", x"0d662fb3", x"1e4abaa3", x"233c6c47", x"1ecbcf17", x"04a400fd", x"f6da4000", x"ae300000", x"63490000", x"6c507359", x"8aa527ae", x"08da66c2", x"dd7cf848"),
	(x"07bd00a4", x"affe8000", x"79430000", x"64c40000", x"2c511448", x"14f26f0d", x"eef9e75e", x"c95e7526", x"a2db00fc", x"87edc000", x"b7cc0000", x"f5920000", x"56db1ea4", x"616f895d", x"24b7214d", x"71f294c0"),
	(x"a03700a9", x"25b60000", x"876e0000", x"79b00000", x"35785be7", x"0d6822ea", x"75d6da86", x"2c533b85", x"803100f9", x"3e66c000", x"36640000", x"30860000", x"8ba26725", x"a263da9f", x"71443c50", x"5121edd1"),
	(x"56b700ac", x"11f5c000", x"a3690000", x"f68d0000", x"144f601c", x"07d0f744", x"b813519f", x"fbc681b4", x"264e00f8", x"4f514000", x"2f980000", x"a65d0000", x"b1290ad8", x"49a9746c", x"5d297bdf", x"fdaf8159"),
	(x"064800a8", x"54818000", x"9e920000", x"ef6b0000", x"0ff3361a", x"e6a28c19", x"59bb9d09", x"80dd570d", x"d0ce00fd", x"7b128000", x"0b9f0000", x"29600000", x"901e3123", x"4311a1c2", x"90ecf0c6", x"2a3a3b68"),
	(x"f0c800ad", x"60c24000", x"ba950000", x"60560000", x"2ec40de1", x"ec1a59b7", x"947e1610", x"5748ed3c", x"76b100fc", x"0a250000", x"12630000", x"bfbb0000", x"aa955cde", x"a8db0f31", x"bc81b749", x"86b457e0"),
	(x"e8870170", x"9d720000", x"12db0000", x"d4220000", x"f2886b27", x"a921e543", x"4ef8b518", x"618813b1", x"b4370060", x"0c4c0000", x"56c20000", x"5cae0000", x"94541f3f", x"3b3ef825", x"1b365f3d", x"f3d45758"),
	(x"1e070175", x"a931c000", x"36dc0000", x"5b1f0000", x"d3bf50dc", x"a39930ed", x"833d3e01", x"b61da980", x"12480061", x"7d7b8000", x"4f3e0000", x"ca750000", x"aedf72c2", x"d0f456d6", x"375b18b2", x"5f5a3bd0"),
	(x"4ef80171", x"ec458000", x"0b270000", x"42f90000", x"c80306da", x"42eb4bb0", x"6295f297", x"cd067f39", x"e4c80064", x"49384000", x"6b390000", x"45480000", x"8fe84939", x"da4c8378", x"fa9e93ab", x"88cf81e1"),
	(x"b8780174", x"d8064000", x"2f200000", x"cdc40000", x"e9343d21", x"48539e1e", x"af50798e", x"1a93c508", x"42b70065", x"380fc000", x"72c50000", x"d3930000", x"b56324c4", x"31862d8b", x"d6f3d424", x"2441ed69"),
	(x"1ff20179", x"524ec000", x"d10d0000", x"d0b00000", x"f01d728e", x"51c9d3f9", x"347f4456", x"ff9e8bab", x"605d0060", x"8184c000", x"f36d0000", x"16870000", x"681a5d45", x"f28a7e49", x"8300c939", x"04929478"),
	(x"e972017c", x"660d0000", x"f50a0000", x"5f8d0000", x"d12a4975", x"5b710657", x"f9bacf4f", x"280b319a", x"c6220061", x"f0b34000", x"ea910000", x"805c0000", x"529130b8", x"1940d0ba", x"af6d8eb6", x"a81cf8f0"),
	(x"b98d0178", x"23794000", x"c8f10000", x"466b0000", x"ca961f73", x"ba037d0a", x"181203d9", x"5310e723", x"30a20064", x"c4f08000", x"ce960000", x"0f610000", x"73a60b43", x"13f80514", x"62a805af", x"7f8942c1"),
	(x"4f0d017d", x"173a8000", x"ecf60000", x"c9560000", x"eba12488", x"b0bba8a4", x"d5d788c0", x"84855d12", x"96dd0065", x"b5c70000", x"d76a0000", x"99ba0000", x"492d66be", x"f832abe7", x"4ec54220", x"d3072e49"),
	(x"3ced0170", x"10bac000", x"b7740000", x"9e0b0000", x"0ec6295d", x"6095632f", x"d6ce231c", x"96ced091", x"97280069", x"4eb80000", x"30bb0000", x"12150000", x"6a8f44ec", x"0a6248f3", x"f9873877", x"9a840c62"),
	(x"ca6d0175", x"24f90000", x"93730000", x"11360000", x"2ff112a6", x"6a2db681", x"1b0ba805", x"415b6aa0", x"31570068", x"3f8f8000", x"29470000", x"84ce0000", x"50042911", x"e1a8e600", x"d5ea7ff8", x"360a60ea"),
	(x"9a920171", x"618d4000", x"ae880000", x"08d00000", x"344d44a0", x"8b5fcddc", x"faa36493", x"3a40bc19", x"c7d7006d", x"0bcc4000", x"0d400000", x"0bf30000", x"713312ea", x"eb1033ae", x"182ff4e1", x"e19fdadb"),
	(x"6c120174", x"55ce8000", x"8a8f0000", x"87ed0000", x"157a7f5b", x"81e71872", x"3766ef8a", x"edd50628", x"61a8006c", x"7afbc000", x"14bc0000", x"9d280000", x"4bb87f17", x"00da9d5d", x"3442b36e", x"4d11b653"),
	(x"cb980179", x"df860000", x"74a20000", x"9a990000", x"0c5330f4", x"987d5595", x"ac49d252", x"08d8488b", x"43420069", x"c370c000", x"95140000", x"583c0000", x"96c10696", x"c3d6ce9f", x"61b1ae73", x"6dc2cf42"),
	(x"3d18017c", x"ebc5c000", x"50a50000", x"15a40000", x"2d640b0f", x"92c5803b", x"618c594b", x"df4df2ba", x"e53d0068", x"b2474000", x"8ce80000", x"cee70000", x"ac4a6b6b", x"281c606c", x"4ddce9fc", x"c14ca3ca"),
	(x"6de70178", x"aeb18000", x"6d5e0000", x"0c420000", x"36d85d09", x"73b7fb66", x"802495dd", x"a4562403", x"13bd006d", x"86048000", x"a8ef0000", x"41da0000", x"8d7d5090", x"22a4b5c2", x"801962e5", x"16d919fb"),
	(x"9b67017d", x"9af24000", x"49590000", x"837f0000", x"17ef66f2", x"790f2ec8", x"4de11ec4", x"73c39e32", x"b5c2006c", x"f7330000", x"b1130000", x"d7010000", x"b7f63d6d", x"c96e1b31", x"ac74256a", x"ba577573"),
	(x"9fc30180", x"6c280000", x"e7690000", x"e0360000", x"7bbf15ab", x"f3aa0966", x"453b7806", x"aebf667a", x"405b0030", x"9a540000", x"42670000", x"5fb10000", x"d6c06187", x"5d81863c", x"87922fef", x"79e0422c"),
	(x"69430185", x"586bc000", x"c36e0000", x"6f0b0000", x"5a882e50", x"f912dcc8", x"88fef31f", x"792adc4b", x"e6240031", x"eb638000", x"5b9b0000", x"c96a0000", x"ec4b0c7a", x"b64b28cf", x"abff6860", x"d56e2ea4"),
	(x"39bc0181", x"1d1f8000", x"fe950000", x"76ed0000", x"41347856", x"1860a795", x"69563f89", x"02310af2", x"10a40034", x"df204000", x"7f9c0000", x"46570000", x"cd7c3781", x"bcf3fd61", x"663ae379", x"02fb9495"),
	(x"cf3c0184", x"295c4000", x"da920000", x"f9d00000", x"600343ad", x"12d8723b", x"a493b490", x"d5a4b0c3", x"b6db0035", x"ae17c000", x"66600000", x"d08c0000", x"f7f75a7c", x"57395392", x"4a57a4f6", x"ae75f81d"),
	(x"68b60189", x"a314c000", x"24bf0000", x"e4a40000", x"792a0c02", x"0b423fdc", x"3fbc8948", x"30a9fe60", x"94310030", x"179cc000", x"e7c80000", x"15980000", x"2a8e23fd", x"94350050", x"1fa4b9eb", x"8ea6810c"),
	(x"9e36018c", x"97570000", x"00b80000", x"6b990000", x"581d37f9", x"01faea72", x"f2790251", x"e73c4451", x"324e0031", x"66ab4000", x"fe340000", x"83430000", x"10054e00", x"7fffaea3", x"33c9fe64", x"2228ed84"),
	(x"cec90188", x"d2234000", x"3d430000", x"727f0000", x"43a161ff", x"e088912f", x"13d1cec7", x"9c2792e8", x"c4ce0034", x"52e88000", x"da330000", x"0c7e0000", x"313275fb", x"75477b0d", x"fe0c757d", x"f5bd57b5"),
	(x"3849018d", x"e6608000", x"19440000", x"fd420000", x"62965a04", x"ea304481", x"de1445de", x"4bb228d9", x"62b10035", x"23df0000", x"c3cf0000", x"9aa50000", x"0bb91806", x"9e8dd5fe", x"d26132f2", x"59333b3d"),
	(x"4ba90180", x"e1e0c000", x"42c60000", x"aa1f0000", x"87f157d1", x"3a1e8f0a", x"dd0dee02", x"59f9a55a", x"63440039", x"d8a00000", x"241e0000", x"110a0000", x"281b3a54", x"6cdd36ea", x"652348a5", x"10b01916"),
	(x"bd290185", x"d5a30000", x"66c10000", x"25220000", x"a6c66c2a", x"30a65aa4", x"10c8651b", x"8e6c1f6b", x"c53b0038", x"a9978000", x"3de20000", x"87d10000", x"129057a9", x"87179819", x"494e0f2a", x"bc3e759e"),
	(x"edd60181", x"90d74000", x"5b3a0000", x"3cc40000", x"bd7a3a2c", x"d1d421f9", x"f160a98d", x"f577c9d2", x"33bb003d", x"9dd44000", x"19e50000", x"08ec0000", x"33a76c52", x"8daf4db7", x"848b8433", x"6babcfaf"),
	(x"1b560184", x"a4948000", x"7f3d0000", x"b3f90000", x"9c4d01d7", x"db6cf457", x"3ca52294", x"22e273e3", x"95c4003c", x"ece3c000", x"00190000", x"9e370000", x"092c01af", x"6665e344", x"a8e6c3bc", x"c725a327"),
	(x"bcdc0189", x"2edc0000", x"81100000", x"ae8d0000", x"85644e78", x"c2f6b9b0", x"a78a1f4c", x"c7ef3d40", x"b72e0039", x"5568c000", x"81b10000", x"5b230000", x"d455782e", x"a569b086", x"fd15dea1", x"e7f6da36"),
	(x"4a5c018c", x"1a9fc000", x"a5170000", x"21b00000", x"a4537583", x"c84e6c1e", x"6a4f9455", x"107a8771", x"11510038", x"245f4000", x"984d0000", x"cdf80000", x"eede15d3", x"4ea31e75", x"d178992e", x"4b78b6be"),
	(x"1aa30188", x"5feb8000", x"98ec0000", x"38560000", x"bfef2385", x"293c1743", x"8be758c3", x"6b6151c8", x"e7d1003d", x"101c8000", x"bc4a0000", x"42c50000", x"cfe92e28", x"441bcbdb", x"1cbd1237", x"9ced0c8f"),
	(x"ec23018d", x"6ba84000", x"bceb0000", x"b76b0000", x"9ed8187e", x"2384c2ed", x"4622d3da", x"bcf4ebf9", x"41ae003c", x"612b0000", x"a5b60000", x"d41e0000", x"f56243d5", x"afd16528", x"30d055b8", x"30636007"),
	(x"1ceb0120", x"0b6a0000", x"067e0000", x"d73d0000", x"b01c159f", x"cf9e9b5a", x"d25cc5ca", x"ebbc06c5", x"371f00c0", x"6b0e0000", x"b7d50000", x"6ba50000", x"5ff71f0b", x"070a6a19", x"8c51e2f1", x"b6d737e7"),
	(x"ea6b0125", x"3f29c000", x"22790000", x"58000000", x"912b2e64", x"c5264ef4", x"1f994ed3", x"3c29bcf4", x"916000c1", x"1a398000", x"ae290000", x"fd7e0000", x"657c72f6", x"ecc0c4ea", x"a03ca57e", x"1a595b6f"),
	(x"ba940121", x"7a5d8000", x"1f820000", x"41e60000", x"8a977862", x"245435a9", x"fe318245", x"47326a4d", x"67e000c4", x"2e7a4000", x"8a2e0000", x"72430000", x"444b490d", x"e6781144", x"6df92e67", x"cdcce15e"),
	(x"4c140124", x"4e1e4000", x"3b850000", x"cedb0000", x"aba04399", x"2eece007", x"33f4095c", x"90a7d07c", x"c19f00c5", x"5f4dc000", x"93d20000", x"e4980000", x"7ec024f0", x"0db2bfb7", x"419469e8", x"61428dd6"),
	(x"eb9e0129", x"c456c000", x"c5a80000", x"d3af0000", x"b2890c36", x"3776ade0", x"a8db3484", x"75aa9edf", x"e37500c0", x"e6c6c000", x"127a0000", x"218c0000", x"a3b95d71", x"cebeec75", x"146774f5", x"4191f4c7"),
	(x"1d1e012c", x"f0150000", x"e1af0000", x"5c920000", x"93be37cd", x"3dce784e", x"651ebf9d", x"a23f24ee", x"450a00c1", x"97f14000", x"0b860000", x"b7570000", x"9932308c", x"25744286", x"380a337a", x"ed1f984f"),
	(x"4de10128", x"b5614000", x"dc540000", x"45740000", x"880261cb", x"dcbc0313", x"84b6730b", x"d924f257", x"b38a00c4", x"a3b28000", x"2f810000", x"386a0000", x"b8050b77", x"2fcc9728", x"f5cfb863", x"3a8a227e"),
	(x"bb61012d", x"81228000", x"f8530000", x"ca490000", x"a9355a30", x"d604d6bd", x"4973f812", x"0eb14866", x"15f500c5", x"d2850000", x"367d0000", x"aeb10000", x"828e668a", x"c40639db", x"d9a2ffec", x"96044ef6"),
	(x"c8810120", x"86a2c000", x"a3d10000", x"9d140000", x"4c5257e5", x"062a1d36", x"4a6a53ce", x"1cfac5e5", x"140000c9", x"29fa0000", x"d1ac0000", x"251e0000", x"a12c44d8", x"3656dacf", x"6ee085bb", x"df876cdd"),
	(x"3e010125", x"b2e10000", x"87d60000", x"12290000", x"6d656c1e", x"0c92c898", x"87afd8d7", x"cb6f7fd4", x"b27f00c8", x"58cd8000", x"c8500000", x"b3c50000", x"9ba72925", x"dd9c743c", x"428dc234", x"73090055"),
	(x"6efe0121", x"f7954000", x"ba2d0000", x"0bcf0000", x"76d93a18", x"ede0b3c5", x"66071441", x"b074a96d", x"44ff00cd", x"6c8e4000", x"ec570000", x"3cf80000", x"ba9012de", x"d724a192", x"8f48492d", x"a49cba64"),
	(x"987e0124", x"c3d68000", x"9e2a0000", x"84f20000", x"57ee01e3", x"e758666b", x"abc29f58", x"67e1135c", x"e28000cc", x"1db9c000", x"f5ab0000", x"aa230000", x"801b7f23", x"3cee0f61", x"a3250ea2", x"0812d6ec"),
	(x"3ff40129", x"499e0000", x"60070000", x"99860000", x"4ec74e4c", x"fec22b8c", x"30eda280", x"82ec5dff", x"c06a00c9", x"a432c000", x"74030000", x"6f370000", x"5d6206a2", x"ffe25ca3", x"f6d613bf", x"28c1affd"),
	(x"c974012c", x"7dddc000", x"44000000", x"16bb0000", x"6ff075b7", x"f47afe22", x"fd282999", x"5579e7ce", x"661500c8", x"d5054000", x"6dff0000", x"f9ec0000", x"67e96b5f", x"1428f250", x"dabb5430", x"844fc375"),
	(x"998b0128", x"38a98000", x"79fb0000", x"0f5d0000", x"744c23b1", x"1508857f", x"1c80e50f", x"2e623177", x"909500cd", x"e1468000", x"49f80000", x"76d10000", x"46de50a4", x"1e9027fe", x"177edf29", x"53da7944"),
	(x"6f0b012d", x"0cea4000", x"5dfc0000", x"80600000", x"557b184a", x"1fb050d1", x"d1456e16", x"f9f78b46", x"36ea00cc", x"90710000", x"50040000", x"e00a0000", x"7c553d59", x"f55a890d", x"3b1398a6", x"ff5415cc"),
	(x"6baf01d0", x"fa300000", x"f3cc0000", x"e3290000", x"392b6b13", x"9515777f", x"d99f08d4", x"248b730e", x"c3730090", x"fd160000", x"a3700000", x"68ba0000", x"1d6361b3", x"61b51400", x"10f59223", x"3ce32293"),
	(x"9d2f01d5", x"ce73c000", x"d7cb0000", x"6c140000", x"181c50e8", x"9fada2d1", x"145a83cd", x"f31ec93f", x"650c0091", x"8c218000", x"ba8c0000", x"fe610000", x"27e80c4e", x"8a7fbaf3", x"3c98d5ac", x"906d4e1b"),
	(x"cdd001d1", x"8b078000", x"ea300000", x"75f20000", x"03a006ee", x"7edfd98c", x"f5f24f5b", x"88051f86", x"938c0094", x"b8624000", x"9e8b0000", x"715c0000", x"06df37b5", x"80c76f5d", x"f15d5eb5", x"47f8f42a"),
	(x"3b5001d4", x"bf444000", x"ce370000", x"facf0000", x"22973d15", x"74670c22", x"3837c442", x"5f90a5b7", x"35f30095", x"c955c000", x"87770000", x"e7870000", x"3c545a48", x"6b0dc1ae", x"dd30193a", x"eb7698a2"),
	(x"9cda01d9", x"350cc000", x"301a0000", x"e7bb0000", x"3bbe72ba", x"6dfd41c5", x"a318f99a", x"ba9deb14", x"17190090", x"70dec000", x"06df0000", x"22930000", x"e12d23c9", x"a801926c", x"88c30427", x"cba5e1b3"),
	(x"6a5a01dc", x"014f0000", x"141d0000", x"68860000", x"1a894941", x"6745946b", x"6edd7283", x"6d085125", x"b1660091", x"01e94000", x"1f230000", x"b4480000", x"dba64e34", x"43cb3c9f", x"a4ae43a8", x"672b8d3b"),
	(x"3aa501d8", x"443b4000", x"29e60000", x"71600000", x"01351f47", x"8637ef36", x"8f75be15", x"1613879c", x"47e60094", x"35aa8000", x"3b240000", x"3b750000", x"fa9175cf", x"4973e931", x"696bc8b1", x"b0be370a"),
	(x"cc2501dd", x"70788000", x"0de10000", x"fe5d0000", x"200224bc", x"8c8f3a98", x"42b0350c", x"c1863dad", x"e1990095", x"449d0000", x"22d80000", x"adae0000", x"c01a1832", x"a2b947c2", x"45068f3e", x"1c305b82"),
	(x"bfc501d0", x"77f8c000", x"56630000", x"a9000000", x"c5652969", x"5ca1f113", x"41a99ed0", x"d3cdb02e", x"e06c0099", x"bfe20000", x"c5090000", x"26010000", x"e3b83a60", x"50e9a4d6", x"f244f569", x"55b379a9"),
	(x"494501d5", x"43bb0000", x"72640000", x"263d0000", x"e4521292", x"561924bd", x"8c6c15c9", x"04580a1f", x"46130098", x"ced58000", x"dcf50000", x"b0da0000", x"d933579d", x"bb230a25", x"de29b2e6", x"f93d1521"),
	(x"19ba01d1", x"06cf4000", x"4f9f0000", x"3fdb0000", x"ffee4494", x"b76b5fe0", x"6dc4d95f", x"7f43dca6", x"b093009d", x"fa964000", x"f8f20000", x"3fe70000", x"f8046c66", x"b19bdf8b", x"13ec39ff", x"2ea8af10"),
	(x"ef3a01d4", x"328c8000", x"6b980000", x"b0e60000", x"ded97f6f", x"bdd38a4e", x"a0015246", x"a8d66697", x"16ec009c", x"8ba1c000", x"e10e0000", x"a93c0000", x"c28f019b", x"5a517178", x"3f817e70", x"8226c398"),
	(x"48b001d9", x"b8c40000", x"95b50000", x"ad920000", x"c7f030c0", x"a449c7a9", x"3b2e6f9e", x"4ddb2834", x"34060099", x"322ac000", x"60a60000", x"6c280000", x"1ff6781a", x"995d22ba", x"6a72636d", x"a2f5ba89"),
	(x"be3001dc", x"8c87c000", x"b1b20000", x"22af0000", x"e6c70b3b", x"aef11207", x"f6ebe487", x"9a4e9205", x"92790098", x"431d4000", x"795a0000", x"faf30000", x"257d15e7", x"72978c49", x"461f24e2", x"0e7bd601"),
	(x"eecf01d8", x"c9f38000", x"8c490000", x"3b490000", x"fd7b5d3d", x"4f83695a", x"17432811", x"e15544bc", x"64f9009d", x"775e8000", x"5d5d0000", x"75ce0000", x"044a2e1c", x"782f59e7", x"8bdaaffb", x"d9ee6c30"),
	(x"184f01dd", x"fdb04000", x"a84e0000", x"b4740000", x"dc4c66c6", x"453bbcf4", x"da86a308", x"36c0fe8d", x"c286009c", x"06690000", x"44a10000", x"e3150000", x"3ec143e1", x"93e5f714", x"a7b7e874", x"756000b8"),
	(x"b4370060", x"0c4c0000", x"56c20000", x"5cae0000", x"94541f3f", x"3b3ef825", x"1b365f3d", x"f3d45758", x"5cb00110", x"913e0000", x"44190000", x"888c0000", x"66dc7418", x"921f1d66", x"55ceea25", x"925c44e9"),
	(x"42b70065", x"380fc000", x"72c50000", x"d3930000", x"b56324c4", x"31862d8b", x"d6f3d424", x"2441ed69", x"facf0111", x"e0098000", x"5de50000", x"1e570000", x"5c5719e5", x"79d5b395", x"79a3adaa", x"3ed22861"),
	(x"12480061", x"7d7b8000", x"4f3e0000", x"ca750000", x"aedf72c2", x"d0f456d6", x"375b18b2", x"5f5a3bd0", x"0c4f0114", x"d44a4000", x"79e20000", x"916a0000", x"7d60221e", x"736d663b", x"b46626b3", x"e9479250"),
	(x"e4c80064", x"49384000", x"6b390000", x"45480000", x"8fe84939", x"da4c8378", x"fa9e93ab", x"88cf81e1", x"aa300115", x"a57dc000", x"601e0000", x"07b10000", x"47eb4fe3", x"98a7c8c8", x"980b613c", x"45c9fed8"),
	(x"43420069", x"c370c000", x"95140000", x"583c0000", x"96c10696", x"c3d6ce9f", x"61b1ae73", x"6dc2cf42", x"88da0110", x"1cf6c000", x"e1b60000", x"c2a50000", x"9a923662", x"5bab9b0a", x"cdf87c21", x"651a87c9"),
	(x"b5c2006c", x"f7330000", x"b1130000", x"d7010000", x"b7f63d6d", x"c96e1b31", x"ac74256a", x"ba577573", x"2ea50111", x"6dc14000", x"f84a0000", x"547e0000", x"a0195b9f", x"b06135f9", x"e1953bae", x"c994eb41"),
	(x"e53d0068", x"b2474000", x"8ce80000", x"cee70000", x"ac4a6b6b", x"281c606c", x"4ddce9fc", x"c14ca3ca", x"d8250114", x"59828000", x"dc4d0000", x"db430000", x"812e6064", x"bad9e057", x"2c50b0b7", x"1e015170"),
	(x"13bd006d", x"86048000", x"a8ef0000", x"41da0000", x"8d7d5090", x"22a4b5c2", x"801962e5", x"16d919fb", x"7e5a0115", x"28b50000", x"c5b10000", x"4d980000", x"bba50d99", x"51134ea4", x"003df738", x"b28f3df8"),
	(x"605d0060", x"8184c000", x"f36d0000", x"16870000", x"681a5d45", x"f28a7e49", x"8300c939", x"04929478", x"7faf0119", x"d3ca0000", x"22600000", x"c6370000", x"98072fcb", x"a343adb0", x"b77f8d6f", x"fb0c1fd3"),
	(x"96dd0065", x"b5c70000", x"d76a0000", x"99ba0000", x"492d66be", x"f832abe7", x"4ec54220", x"d3072e49", x"d9d00118", x"a2fd8000", x"3b9c0000", x"50ec0000", x"a28c4236", x"48890343", x"9b12cae0", x"5782735b"),
	(x"c6220061", x"f0b34000", x"ea910000", x"805c0000", x"529130b8", x"1940d0ba", x"af6d8eb6", x"a81cf8f0", x"2f50011d", x"96be4000", x"1f9b0000", x"dfd10000", x"83bb79cd", x"4231d6ed", x"56d741f9", x"8017c96a"),
	(x"30a20064", x"c4f08000", x"ce960000", x"0f610000", x"73a60b43", x"13f80514", x"62a805af", x"7f8942c1", x"892f011c", x"e789c000", x"06670000", x"490a0000", x"b9301430", x"a9fb781e", x"7aba0676", x"2c99a5e2"),
	(x"97280069", x"4eb80000", x"30bb0000", x"12150000", x"6a8f44ec", x"0a6248f3", x"f9873877", x"9a840c62", x"abc50119", x"5e02c000", x"87cf0000", x"8c1e0000", x"64496db1", x"6af72bdc", x"2f491b6b", x"0c4adcf3"),
	(x"61a8006c", x"7afbc000", x"14bc0000", x"9d280000", x"4bb87f17", x"00da9d5d", x"3442b36e", x"4d11b653", x"0dba0118", x"2f354000", x"9e330000", x"1ac50000", x"5ec2004c", x"813d852f", x"03245ce4", x"a0c4b07b"),
	(x"31570068", x"3f8f8000", x"29470000", x"84ce0000", x"50042911", x"e1a8e600", x"d5ea7ff8", x"360a60ea", x"fb3a011d", x"1b768000", x"ba340000", x"95f80000", x"7ff53bb7", x"8b855081", x"cee1d7fd", x"77510a4a"),
	(x"c7d7006d", x"0bcc4000", x"0d400000", x"0bf30000", x"713312ea", x"eb1033ae", x"182ff4e1", x"e19fdadb", x"5d45011c", x"6a410000", x"a3c80000", x"03230000", x"457e564a", x"604ffe72", x"e28c9072", x"dbdf66c2"),
	(x"c3730090", x"fd160000", x"a3700000", x"68ba0000", x"1d6361b3", x"61b51400", x"10f59223", x"3ce32293", x"a8dc0140", x"07260000", x"50bc0000", x"8b930000", x"24480aa0", x"f4a0637f", x"c96a9af7", x"1868519d"),
	(x"35f30095", x"c955c000", x"87770000", x"e7870000", x"3c545a48", x"6b0dc1ae", x"dd30193a", x"eb7698a2", x"0ea30141", x"76118000", x"49400000", x"1d480000", x"1ec3675d", x"1f6acd8c", x"e507dd78", x"b4e63d15"),
	(x"650c0091", x"8c218000", x"ba8c0000", x"fe610000", x"27e80c4e", x"8a7fbaf3", x"3c98d5ac", x"906d4e1b", x"f8230144", x"42524000", x"6d470000", x"92750000", x"3ff45ca6", x"15d21822", x"28c25661", x"63738724"),
	(x"938c0094", x"b8624000", x"9e8b0000", x"715c0000", x"06df37b5", x"80c76f5d", x"f15d5eb5", x"47f8f42a", x"5e5c0145", x"3365c000", x"74bb0000", x"04ae0000", x"057f315b", x"fe18b6d1", x"04af11ee", x"cffdebac"),
	(x"34060099", x"322ac000", x"60a60000", x"6c280000", x"1ff6781a", x"995d22ba", x"6a72636d", x"a2f5ba89", x"7cb60140", x"8aeec000", x"f5130000", x"c1ba0000", x"d80648da", x"3d14e513", x"515c0cf3", x"ef2e92bd"),
	(x"c286009c", x"06690000", x"44a10000", x"e3150000", x"3ec143e1", x"93e5f714", x"a7b7e874", x"756000b8", x"dac90141", x"fbd94000", x"ecef0000", x"57610000", x"e28d2527", x"d6de4be0", x"7d314b7c", x"43a0fe35"),
	(x"92790098", x"431d4000", x"795a0000", x"faf30000", x"257d15e7", x"72978c49", x"461f24e2", x"0e7bd601", x"2c490144", x"cf9a8000", x"c8e80000", x"d85c0000", x"c3ba1edc", x"dc669e4e", x"b0f4c065", x"94354404"),
	(x"64f9009d", x"775e8000", x"5d5d0000", x"75ce0000", x"044a2e1c", x"782f59e7", x"8bdaaffb", x"d9ee6c30", x"8a360145", x"bead0000", x"d1140000", x"4e870000", x"f9317321", x"37ac30bd", x"9c9987ea", x"38bb288c"),
	(x"17190090", x"70dec000", x"06df0000", x"22930000", x"e12d23c9", x"a801926c", x"88c30427", x"cba5e1b3", x"8bc30149", x"45d20000", x"36c50000", x"c5280000", x"da935173", x"c5fcd3a9", x"2bdbfdbd", x"71380aa7"),
	(x"e1990095", x"449d0000", x"22d80000", x"adae0000", x"c01a1832", x"a2b947c2", x"45068f3e", x"1c305b82", x"2dbc0148", x"34e58000", x"2f390000", x"53f30000", x"e0183c8e", x"2e367d5a", x"07b6ba32", x"ddb6662f"),
	(x"b1660091", x"01e94000", x"1f230000", x"b4480000", x"dba64e34", x"43cb3c9f", x"a4ae43a8", x"672b8d3b", x"db3c014d", x"00a64000", x"0b3e0000", x"dcce0000", x"c12f0775", x"248ea8f4", x"ca73312b", x"0a23dc1e"),
	(x"47e60094", x"35aa8000", x"3b240000", x"3b750000", x"fa9175cf", x"4973e931", x"696bc8b1", x"b0be370a", x"7d43014c", x"7191c000", x"12c20000", x"4a150000", x"fba46a88", x"cf440607", x"e61e76a4", x"a6adb096"),
	(x"e06c0099", x"bfe20000", x"c5090000", x"26010000", x"e3b83a60", x"50e9a4d6", x"f244f569", x"55b379a9", x"5fa90149", x"c81ac000", x"936a0000", x"8f010000", x"26dd1309", x"0c4855c5", x"b3ed6bb9", x"867ec987"),
	(x"16ec009c", x"8ba1c000", x"e10e0000", x"a93c0000", x"c28f019b", x"5a517178", x"3f817e70", x"8226c398", x"f9d60148", x"b92d4000", x"8a960000", x"19da0000", x"1c567ef4", x"e782fb36", x"9f802c36", x"2af0a50f"),
	(x"46130098", x"ced58000", x"dcf50000", x"b0da0000", x"d933579d", x"bb230a25", x"de29b2e6", x"f93d1521", x"0f56014d", x"8d6e8000", x"ae910000", x"96e70000", x"3d61450f", x"ed3a2e98", x"5245a72f", x"fd651f3e"),
	(x"b093009d", x"fa964000", x"f8f20000", x"3fe70000", x"f8046c66", x"b19bdf8b", x"13ec39ff", x"2ea8af10", x"a929014c", x"fc590000", x"b76d0000", x"003c0000", x"07ea28f2", x"06f0806b", x"7e28e0a0", x"51eb73b6"),
	(x"405b0030", x"9a540000", x"42670000", x"5fb10000", x"d6c06187", x"5d81863c", x"87922fef", x"79e0422c", x"df9801b0", x"f67c0000", x"a50e0000", x"bf870000", x"ad7f742c", x"ae2b8f5a", x"c2a957e9", x"d75f2456"),
	(x"b6db0035", x"ae17c000", x"66600000", x"d08c0000", x"f7f75a7c", x"57395392", x"4a57a4f6", x"ae75f81d", x"79e701b1", x"874b8000", x"bcf20000", x"295c0000", x"97f419d1", x"45e121a9", x"eec41066", x"7bd148de"),
	(x"e6240031", x"eb638000", x"5b9b0000", x"c96a0000", x"ec4b0c7a", x"b64b28cf", x"abff6860", x"d56e2ea4", x"8f6701b4", x"b3084000", x"98f50000", x"a6610000", x"b6c3222a", x"4f59f407", x"23019b7f", x"ac44f2ef"),
	(x"10a40034", x"df204000", x"7f9c0000", x"46570000", x"cd7c3781", x"bcf3fd61", x"663ae379", x"02fb9495", x"291801b5", x"c23fc000", x"81090000", x"30ba0000", x"8c484fd7", x"a4935af4", x"0f6cdcf0", x"00ca9e67"),
	(x"b72e0039", x"5568c000", x"81b10000", x"5b230000", x"d455782e", x"a569b086", x"fd15dea1", x"e7f6da36", x"0bf201b0", x"7bb4c000", x"00a10000", x"f5ae0000", x"51313656", x"679f0936", x"5a9fc1ed", x"2019e776"),
	(x"41ae003c", x"612b0000", x"a5b60000", x"d41e0000", x"f56243d5", x"afd16528", x"30d055b8", x"30636007", x"ad8d01b1", x"0a834000", x"195d0000", x"63750000", x"6bba5bab", x"8c55a7c5", x"76f28662", x"8c978bfe"),
	(x"11510038", x"245f4000", x"984d0000", x"cdf80000", x"eede15d3", x"4ea31e75", x"d178992e", x"4b78b6be", x"5b0d01b4", x"3ec08000", x"3d5a0000", x"ec480000", x"4a8d6050", x"86ed726b", x"bb370d7b", x"5b0231cf"),
	(x"e7d1003d", x"101c8000", x"bc4a0000", x"42c50000", x"cfe92e28", x"441bcbdb", x"1cbd1237", x"9ced0c8f", x"fd7201b5", x"4ff70000", x"24a60000", x"7a930000", x"70060dad", x"6d27dc98", x"975a4af4", x"f78c5d47"),
	(x"94310030", x"179cc000", x"e7c80000", x"15980000", x"2a8e23fd", x"94350050", x"1fa4b9eb", x"8ea6810c", x"fc8701b9", x"b4880000", x"c3770000", x"f13c0000", x"53a42fff", x"9f773f8c", x"201830a3", x"be0f7f6c"),
	(x"62b10035", x"23df0000", x"c3cf0000", x"9aa50000", x"0bb91806", x"9e8dd5fe", x"d26132f2", x"59333b3d", x"5af801b8", x"c5bf8000", x"da8b0000", x"67e70000", x"692f4202", x"74bd917f", x"0c75772c", x"128113e4"),
	(x"324e0031", x"66ab4000", x"fe340000", x"83430000", x"10054e00", x"7fffaea3", x"33c9fe64", x"2228ed84", x"ac7801bd", x"f1fc4000", x"fe8c0000", x"e8da0000", x"481879f9", x"7e0544d1", x"c1b0fc35", x"c514a9d5"),
	(x"c4ce0034", x"52e88000", x"da330000", x"0c7e0000", x"313275fb", x"75477b0d", x"fe0c757d", x"f5bd57b5", x"0a0701bc", x"80cbc000", x"e7700000", x"7e010000", x"72931404", x"95cfea22", x"edddbbba", x"699ac55d"),
	(x"63440039", x"d8a00000", x"241e0000", x"110a0000", x"281b3a54", x"6cdd36ea", x"652348a5", x"10b01916", x"28ed01b9", x"3940c000", x"66d80000", x"bb150000", x"afea6d85", x"56c3b9e0", x"b82ea6a7", x"4949bc4c"),
	(x"95c4003c", x"ece3c000", x"00190000", x"9e370000", x"092c01af", x"6665e344", x"a8e6c3bc", x"c725a327", x"8e9201b8", x"48774000", x"7f240000", x"2dce0000", x"95610078", x"bd091713", x"9443e128", x"e5c7d0c4"),
	(x"c53b0038", x"a9978000", x"3de20000", x"87d10000", x"129057a9", x"87179819", x"494e0f2a", x"bc3e759e", x"781201bd", x"7c348000", x"5b230000", x"a2f30000", x"b4563b83", x"b7b1c2bd", x"59866a31", x"32526af5"),
	(x"33bb003d", x"9dd44000", x"19e50000", x"08ec0000", x"33a76c52", x"8daf4db7", x"848b8433", x"6babcfaf", x"de6d01bc", x"0d030000", x"42df0000", x"34280000", x"8edd567e", x"5c7b6c4e", x"75eb2dbe", x"9edc067d"),
	(x"371f00c0", x"6b0e0000", x"b7d50000", x"6ba50000", x"5ff71f0b", x"070a6a19", x"8c51e2f1", x"b6d737e7", x"2bf401e0", x"60640000", x"b1ab0000", x"bc980000", x"efeb0a94", x"c894f143", x"5e0d273b", x"5d6b3122"),
	(x"c19f00c5", x"5f4dc000", x"93d20000", x"e4980000", x"7ec024f0", x"0db2bfb7", x"419469e8", x"61428dd6", x"8d8b01e1", x"11538000", x"a8570000", x"2a430000", x"d5606769", x"235e5fb0", x"726060b4", x"f1e55daa"),
	(x"916000c1", x"1a398000", x"ae290000", x"fd7e0000", x"657c72f6", x"ecc0c4ea", x"a03ca57e", x"1a595b6f", x"7b0b01e4", x"25104000", x"8c500000", x"a57e0000", x"f4575c92", x"29e68a1e", x"bfa5ebad", x"2670e79b"),
	(x"67e000c4", x"2e7a4000", x"8a2e0000", x"72430000", x"444b490d", x"e6781144", x"6df92e67", x"cdcce15e", x"dd7401e5", x"5427c000", x"95ac0000", x"33a50000", x"cedc316f", x"c22c24ed", x"93c8ac22", x"8afe8b13"),
	(x"c06a00c9", x"a432c000", x"74030000", x"6f370000", x"5d6206a2", x"ffe25ca3", x"f6d613bf", x"28c1affd", x"ff9e01e0", x"edacc000", x"14040000", x"f6b10000", x"13a548ee", x"0120772f", x"c63bb13f", x"aa2df202"),
	(x"36ea00cc", x"90710000", x"50040000", x"e00a0000", x"7c553d59", x"f55a890d", x"3b1398a6", x"ff5415cc", x"59e101e1", x"9c9b4000", x"0df80000", x"606a0000", x"292e2513", x"eaead9dc", x"ea56f6b0", x"06a39e8a"),
	(x"661500c8", x"d5054000", x"6dff0000", x"f9ec0000", x"67e96b5f", x"1428f250", x"dabb5430", x"844fc375", x"af6101e4", x"a8d88000", x"29ff0000", x"ef570000", x"08191ee8", x"e0520c72", x"27937da9", x"d13624bb"),
	(x"909500cd", x"e1468000", x"49f80000", x"76d10000", x"46de50a4", x"1e9027fe", x"177edf29", x"53da7944", x"091e01e5", x"d9ef0000", x"30030000", x"798c0000", x"32927315", x"0b98a281", x"0bfe3a26", x"7db84833"),
	(x"e37500c0", x"e6c6c000", x"127a0000", x"218c0000", x"a3b95d71", x"cebeec75", x"146774f5", x"4191f4c7", x"08eb01e9", x"22900000", x"d7d20000", x"f2230000", x"11305147", x"f9c84195", x"bcbc4071", x"343b6a18"),
	(x"15f500c5", x"d2850000", x"367d0000", x"aeb10000", x"828e668a", x"c40639db", x"d9a2ffec", x"96044ef6", x"ae9401e8", x"53a78000", x"ce2e0000", x"64f80000", x"2bbb3cba", x"1202ef66", x"90d107fe", x"98b50690"),
	(x"450a00c1", x"97f14000", x"0b860000", x"b7570000", x"9932308c", x"25744286", x"380a337a", x"ed1f984f", x"581401ed", x"67e44000", x"ea290000", x"ebc50000", x"0a8c0741", x"18ba3ac8", x"5d148ce7", x"4f20bca1"),
	(x"b38a00c4", x"a3b28000", x"2f810000", x"386a0000", x"b8050b77", x"2fcc9728", x"f5cfb863", x"3a8a227e", x"fe6b01ec", x"16d3c000", x"f3d50000", x"7d1e0000", x"30076abc", x"f370943b", x"7179cb68", x"e3aed029"),
	(x"140000c9", x"29fa0000", x"d1ac0000", x"251e0000", x"a12c44d8", x"3656dacf", x"6ee085bb", x"df876cdd", x"dc8101e9", x"af58c000", x"727d0000", x"b80a0000", x"ed7e133d", x"307cc7f9", x"248ad675", x"c37da938"),
	(x"e28000cc", x"1db9c000", x"f5ab0000", x"aa230000", x"801b7f23", x"3cee0f61", x"a3250ea2", x"0812d6ec", x"7afe01e8", x"de6f4000", x"6b810000", x"2ed10000", x"d7f57ec0", x"dbb6690a", x"08e791fa", x"6ff3c5b0"),
	(x"b27f00c8", x"58cd8000", x"c8500000", x"b3c50000", x"9ba72925", x"dd9c743c", x"428dc234", x"73090055", x"8c7e01ed", x"ea2c8000", x"4f860000", x"a1ec0000", x"f6c2453b", x"d10ebca4", x"c5221ae3", x"b8667f81"),
	(x"44ff00cd", x"6c8e4000", x"ec570000", x"3cf80000", x"ba9012de", x"d724a192", x"8f48492d", x"a49cba64", x"2a0101ec", x"9b1b0000", x"567a0000", x"37370000", x"cc4928c6", x"3ac41257", x"e94f5d6c", x"14e81309"),
	(x"5cb00110", x"913e0000", x"44190000", x"888c0000", x"66dc7418", x"921f1d66", x"55ceea25", x"925c44e9", x"e8870170", x"9d720000", x"12db0000", x"d4220000", x"f2886b27", x"a921e543", x"4ef8b518", x"618813b1"),
	(x"aa300115", x"a57dc000", x"601e0000", x"07b10000", x"47eb4fe3", x"98a7c8c8", x"980b613c", x"45c9fed8", x"4ef80171", x"ec458000", x"0b270000", x"42f90000", x"c80306da", x"42eb4bb0", x"6295f297", x"cd067f39"),
	(x"facf0111", x"e0098000", x"5de50000", x"1e570000", x"5c5719e5", x"79d5b395", x"79a3adaa", x"3ed22861", x"b8780174", x"d8064000", x"2f200000", x"cdc40000", x"e9343d21", x"48539e1e", x"af50798e", x"1a93c508"),
	(x"0c4f0114", x"d44a4000", x"79e20000", x"916a0000", x"7d60221e", x"736d663b", x"b46626b3", x"e9479250", x"1e070175", x"a931c000", x"36dc0000", x"5b1f0000", x"d3bf50dc", x"a39930ed", x"833d3e01", x"b61da980"),
	(x"abc50119", x"5e02c000", x"87cf0000", x"8c1e0000", x"64496db1", x"6af72bdc", x"2f491b6b", x"0c4adcf3", x"3ced0170", x"10bac000", x"b7740000", x"9e0b0000", x"0ec6295d", x"6095632f", x"d6ce231c", x"96ced091"),
	(x"5d45011c", x"6a410000", x"a3c80000", x"03230000", x"457e564a", x"604ffe72", x"e28c9072", x"dbdf66c2", x"9a920171", x"618d4000", x"ae880000", x"08d00000", x"344d44a0", x"8b5fcddc", x"faa36493", x"3a40bc19"),
	(x"0dba0118", x"2f354000", x"9e330000", x"1ac50000", x"5ec2004c", x"813d852f", x"03245ce4", x"a0c4b07b", x"6c120174", x"55ce8000", x"8a8f0000", x"87ed0000", x"157a7f5b", x"81e71872", x"3766ef8a", x"edd50628"),
	(x"fb3a011d", x"1b768000", x"ba340000", x"95f80000", x"7ff53bb7", x"8b855081", x"cee1d7fd", x"77510a4a", x"ca6d0175", x"24f90000", x"93730000", x"11360000", x"2ff112a6", x"6a2db681", x"1b0ba805", x"415b6aa0"),
	(x"88da0110", x"1cf6c000", x"e1b60000", x"c2a50000", x"9a923662", x"5bab9b0a", x"cdf87c21", x"651a87c9", x"cb980179", x"df860000", x"74a20000", x"9a990000", x"0c5330f4", x"987d5595", x"ac49d252", x"08d8488b"),
	(x"7e5a0115", x"28b50000", x"c5b10000", x"4d980000", x"bba50d99", x"51134ea4", x"003df738", x"b28f3df8", x"6de70178", x"aeb18000", x"6d5e0000", x"0c420000", x"36d85d09", x"73b7fb66", x"802495dd", x"a4562403"),
	(x"2ea50111", x"6dc14000", x"f84a0000", x"547e0000", x"a0195b9f", x"b06135f9", x"e1953bae", x"c994eb41", x"9b67017d", x"9af24000", x"49590000", x"837f0000", x"17ef66f2", x"790f2ec8", x"4de11ec4", x"73c39e32"),
	(x"d8250114", x"59828000", x"dc4d0000", x"db430000", x"812e6064", x"bad9e057", x"2c50b0b7", x"1e015170", x"3d18017c", x"ebc5c000", x"50a50000", x"15a40000", x"2d640b0f", x"92c5803b", x"618c594b", x"df4df2ba"),
	(x"7faf0119", x"d3ca0000", x"22600000", x"c6370000", x"98072fcb", x"a343adb0", x"b77f8d6f", x"fb0c1fd3", x"1ff20179", x"524ec000", x"d10d0000", x"d0b00000", x"f01d728e", x"51c9d3f9", x"347f4456", x"ff9e8bab"),
	(x"892f011c", x"e789c000", x"06670000", x"490a0000", x"b9301430", x"a9fb781e", x"7aba0676", x"2c99a5e2", x"b98d0178", x"23794000", x"c8f10000", x"466b0000", x"ca961f73", x"ba037d0a", x"181203d9", x"5310e723"),
	(x"d9d00118", x"a2fd8000", x"3b9c0000", x"50ec0000", x"a28c4236", x"48890343", x"9b12cae0", x"5782735b", x"4f0d017d", x"173a8000", x"ecf60000", x"c9560000", x"eba12488", x"b0bba8a4", x"d5d788c0", x"84855d12"),
	(x"2f50011d", x"96be4000", x"1f9b0000", x"dfd10000", x"83bb79cd", x"4231d6ed", x"56d741f9", x"8017c96a", x"e972017c", x"660d0000", x"f50a0000", x"5f8d0000", x"d12a4975", x"5b710657", x"f9bacf4f", x"280b319a"),
	(x"2bf401e0", x"60640000", x"b1ab0000", x"bc980000", x"efeb0a94", x"c894f143", x"5e0d273b", x"5d6b3122", x"1ceb0120", x"0b6a0000", x"067e0000", x"d73d0000", x"b01c159f", x"cf9e9b5a", x"d25cc5ca", x"ebbc06c5"),
	(x"dd7401e5", x"5427c000", x"95ac0000", x"33a50000", x"cedc316f", x"c22c24ed", x"93c8ac22", x"8afe8b13", x"ba940121", x"7a5d8000", x"1f820000", x"41e60000", x"8a977862", x"245435a9", x"fe318245", x"47326a4d"),
	(x"8d8b01e1", x"11538000", x"a8570000", x"2a430000", x"d5606769", x"235e5fb0", x"726060b4", x"f1e55daa", x"4c140124", x"4e1e4000", x"3b850000", x"cedb0000", x"aba04399", x"2eece007", x"33f4095c", x"90a7d07c"),
	(x"7b0b01e4", x"25104000", x"8c500000", x"a57e0000", x"f4575c92", x"29e68a1e", x"bfa5ebad", x"2670e79b", x"ea6b0125", x"3f29c000", x"22790000", x"58000000", x"912b2e64", x"c5264ef4", x"1f994ed3", x"3c29bcf4"),
	(x"dc8101e9", x"af58c000", x"727d0000", x"b80a0000", x"ed7e133d", x"307cc7f9", x"248ad675", x"c37da938", x"c8810120", x"86a2c000", x"a3d10000", x"9d140000", x"4c5257e5", x"062a1d36", x"4a6a53ce", x"1cfac5e5"),
	(x"2a0101ec", x"9b1b0000", x"567a0000", x"37370000", x"cc4928c6", x"3ac41257", x"e94f5d6c", x"14e81309", x"6efe0121", x"f7954000", x"ba2d0000", x"0bcf0000", x"76d93a18", x"ede0b3c5", x"66071441", x"b074a96d"),
	(x"7afe01e8", x"de6f4000", x"6b810000", x"2ed10000", x"d7f57ec0", x"dbb6690a", x"08e791fa", x"6ff3c5b0", x"987e0124", x"c3d68000", x"9e2a0000", x"84f20000", x"57ee01e3", x"e758666b", x"abc29f58", x"67e1135c"),
	(x"8c7e01ed", x"ea2c8000", x"4f860000", x"a1ec0000", x"f6c2453b", x"d10ebca4", x"c5221ae3", x"b8667f81", x"3e010125", x"b2e10000", x"87d60000", x"12290000", x"6d656c1e", x"0c92c898", x"87afd8d7", x"cb6f7fd4"),
	(x"ff9e01e0", x"edacc000", x"14040000", x"f6b10000", x"13a548ee", x"0120772f", x"c63bb13f", x"aa2df202", x"3ff40129", x"499e0000", x"60070000", x"99860000", x"4ec74e4c", x"fec22b8c", x"30eda280", x"82ec5dff"),
	(x"091e01e5", x"d9ef0000", x"30030000", x"798c0000", x"32927315", x"0b98a281", x"0bfe3a26", x"7db84833", x"998b0128", x"38a98000", x"79fb0000", x"0f5d0000", x"744c23b1", x"1508857f", x"1c80e50f", x"2e623177"),
	(x"59e101e1", x"9c9b4000", x"0df80000", x"606a0000", x"292e2513", x"eaead9dc", x"ea56f6b0", x"06a39e8a", x"6f0b012d", x"0cea4000", x"5dfc0000", x"80600000", x"557b184a", x"1fb050d1", x"d1456e16", x"f9f78b46"),
	(x"af6101e4", x"a8d88000", x"29ff0000", x"ef570000", x"08191ee8", x"e0520c72", x"27937da9", x"d13624bb", x"c974012c", x"7dddc000", x"44000000", x"16bb0000", x"6ff075b7", x"f47afe22", x"fd282999", x"5579e7ce"),
	(x"08eb01e9", x"22900000", x"d7d20000", x"f2230000", x"11305147", x"f9c84195", x"bcbc4071", x"343b6a18", x"eb9e0129", x"c456c000", x"c5a80000", x"d3af0000", x"b2890c36", x"3776ade0", x"a8db3484", x"75aa9edf"),
	(x"fe6b01ec", x"16d3c000", x"f3d50000", x"7d1e0000", x"30076abc", x"f370943b", x"7179cb68", x"e3aed029", x"4de10128", x"b5614000", x"dc540000", x"45740000", x"880261cb", x"dcbc0313", x"84b6730b", x"d924f257"),
	(x"ae9401e8", x"53a78000", x"ce2e0000", x"64f80000", x"2bbb3cba", x"1202ef66", x"90d107fe", x"98b50690", x"bb61012d", x"81228000", x"f8530000", x"ca490000", x"a9355a30", x"d604d6bd", x"4973f812", x"0eb14866"),
	(x"581401ed", x"67e44000", x"ea290000", x"ebc50000", x"0a8c0741", x"18ba3ac8", x"5d148ce7", x"4f20bca1", x"1d1e012c", x"f0150000", x"e1af0000", x"5c920000", x"93be37cd", x"3dce784e", x"651ebf9d", x"a23f24ee"),
	(x"a8dc0140", x"07260000", x"50bc0000", x"8b930000", x"24480aa0", x"f4a0637f", x"c96a9af7", x"1868519d", x"6baf01d0", x"fa300000", x"f3cc0000", x"e3290000", x"392b6b13", x"9515777f", x"d99f08d4", x"248b730e"),
	(x"5e5c0145", x"3365c000", x"74bb0000", x"04ae0000", x"057f315b", x"fe18b6d1", x"04af11ee", x"cffdebac", x"cdd001d1", x"8b078000", x"ea300000", x"75f20000", x"03a006ee", x"7edfd98c", x"f5f24f5b", x"88051f86"),
	(x"0ea30141", x"76118000", x"49400000", x"1d480000", x"1ec3675d", x"1f6acd8c", x"e507dd78", x"b4e63d15", x"3b5001d4", x"bf444000", x"ce370000", x"facf0000", x"22973d15", x"74670c22", x"3837c442", x"5f90a5b7"),
	(x"f8230144", x"42524000", x"6d470000", x"92750000", x"3ff45ca6", x"15d21822", x"28c25661", x"63738724", x"9d2f01d5", x"ce73c000", x"d7cb0000", x"6c140000", x"181c50e8", x"9fada2d1", x"145a83cd", x"f31ec93f"),
	(x"5fa90149", x"c81ac000", x"936a0000", x"8f010000", x"26dd1309", x"0c4855c5", x"b3ed6bb9", x"867ec987", x"bfc501d0", x"77f8c000", x"56630000", x"a9000000", x"c5652969", x"5ca1f113", x"41a99ed0", x"d3cdb02e"),
	(x"a929014c", x"fc590000", x"b76d0000", x"003c0000", x"07ea28f2", x"06f0806b", x"7e28e0a0", x"51eb73b6", x"19ba01d1", x"06cf4000", x"4f9f0000", x"3fdb0000", x"ffee4494", x"b76b5fe0", x"6dc4d95f", x"7f43dca6"),
	(x"f9d60148", x"b92d4000", x"8a960000", x"19da0000", x"1c567ef4", x"e782fb36", x"9f802c36", x"2af0a50f", x"ef3a01d4", x"328c8000", x"6b980000", x"b0e60000", x"ded97f6f", x"bdd38a4e", x"a0015246", x"a8d66697"),
	(x"0f56014d", x"8d6e8000", x"ae910000", x"96e70000", x"3d61450f", x"ed3a2e98", x"5245a72f", x"fd651f3e", x"494501d5", x"43bb0000", x"72640000", x"263d0000", x"e4521292", x"561924bd", x"8c6c15c9", x"04580a1f"),
	(x"7cb60140", x"8aeec000", x"f5130000", x"c1ba0000", x"d80648da", x"3d14e513", x"515c0cf3", x"ef2e92bd", x"48b001d9", x"b8c40000", x"95b50000", x"ad920000", x"c7f030c0", x"a449c7a9", x"3b2e6f9e", x"4ddb2834"),
	(x"8a360145", x"bead0000", x"d1140000", x"4e870000", x"f9317321", x"37ac30bd", x"9c9987ea", x"38bb288c", x"eecf01d8", x"c9f38000", x"8c490000", x"3b490000", x"fd7b5d3d", x"4f83695a", x"17432811", x"e15544bc"),
	(x"dac90141", x"fbd94000", x"ecef0000", x"57610000", x"e28d2527", x"d6de4be0", x"7d314b7c", x"43a0fe35", x"184f01dd", x"fdb04000", x"a84e0000", x"b4740000", x"dc4c66c6", x"453bbcf4", x"da86a308", x"36c0fe8d"),
	(x"2c490144", x"cf9a8000", x"c8e80000", x"d85c0000", x"c3ba1edc", x"dc669e4e", x"b0f4c065", x"94354404", x"be3001dc", x"8c87c000", x"b1b20000", x"22af0000", x"e6c70b3b", x"aef11207", x"f6ebe487", x"9a4e9205"),
	(x"8bc30149", x"45d20000", x"36c50000", x"c5280000", x"da935173", x"c5fcd3a9", x"2bdbfdbd", x"71380aa7", x"9cda01d9", x"350cc000", x"301a0000", x"e7bb0000", x"3bbe72ba", x"6dfd41c5", x"a318f99a", x"ba9deb14"),
	(x"7d43014c", x"7191c000", x"12c20000", x"4a150000", x"fba46a88", x"cf440607", x"e61e76a4", x"a6adb096", x"3aa501d8", x"443b4000", x"29e60000", x"71600000", x"01351f47", x"8637ef36", x"8f75be15", x"1613879c"),
	(x"2dbc0148", x"34e58000", x"2f390000", x"53f30000", x"e0183c8e", x"2e367d5a", x"07b6ba32", x"ddb6662f", x"cc2501dd", x"70788000", x"0de10000", x"fe5d0000", x"200224bc", x"8c8f3a98", x"42b0350c", x"c1863dad"),
	(x"db3c014d", x"00a64000", x"0b3e0000", x"dcce0000", x"c12f0775", x"248ea8f4", x"ca73312b", x"0a23dc1e", x"6a5a01dc", x"014f0000", x"141d0000", x"68860000", x"1a894941", x"6745946b", x"6edd7283", x"6d085125"),
	(x"df9801b0", x"f67c0000", x"a50e0000", x"bf870000", x"ad7f742c", x"ae2b8f5a", x"c2a957e9", x"d75f2456", x"9fc30180", x"6c280000", x"e7690000", x"e0360000", x"7bbf15ab", x"f3aa0966", x"453b7806", x"aebf667a"),
	(x"291801b5", x"c23fc000", x"81090000", x"30ba0000", x"8c484fd7", x"a4935af4", x"0f6cdcf0", x"00ca9e67", x"39bc0181", x"1d1f8000", x"fe950000", x"76ed0000", x"41347856", x"1860a795", x"69563f89", x"02310af2"),
	(x"79e701b1", x"874b8000", x"bcf20000", x"295c0000", x"97f419d1", x"45e121a9", x"eec41066", x"7bd148de", x"cf3c0184", x"295c4000", x"da920000", x"f9d00000", x"600343ad", x"12d8723b", x"a493b490", x"d5a4b0c3"),
	(x"8f6701b4", x"b3084000", x"98f50000", x"a6610000", x"b6c3222a", x"4f59f407", x"23019b7f", x"ac44f2ef", x"69430185", x"586bc000", x"c36e0000", x"6f0b0000", x"5a882e50", x"f912dcc8", x"88fef31f", x"792adc4b"),
	(x"28ed01b9", x"3940c000", x"66d80000", x"bb150000", x"afea6d85", x"56c3b9e0", x"b82ea6a7", x"4949bc4c", x"4ba90180", x"e1e0c000", x"42c60000", x"aa1f0000", x"87f157d1", x"3a1e8f0a", x"dd0dee02", x"59f9a55a"),
	(x"de6d01bc", x"0d030000", x"42df0000", x"34280000", x"8edd567e", x"5c7b6c4e", x"75eb2dbe", x"9edc067d", x"edd60181", x"90d74000", x"5b3a0000", x"3cc40000", x"bd7a3a2c", x"d1d421f9", x"f160a98d", x"f577c9d2"),
	(x"8e9201b8", x"48774000", x"7f240000", x"2dce0000", x"95610078", x"bd091713", x"9443e128", x"e5c7d0c4", x"1b560184", x"a4948000", x"7f3d0000", x"b3f90000", x"9c4d01d7", x"db6cf457", x"3ca52294", x"22e273e3"),
	(x"781201bd", x"7c348000", x"5b230000", x"a2f30000", x"b4563b83", x"b7b1c2bd", x"59866a31", x"32526af5", x"bd290185", x"d5a30000", x"66c10000", x"25220000", x"a6c66c2a", x"30a65aa4", x"10c8651b", x"8e6c1f6b"),
	(x"0bf201b0", x"7bb4c000", x"00a10000", x"f5ae0000", x"51313656", x"679f0936", x"5a9fc1ed", x"2019e776", x"bcdc0189", x"2edc0000", x"81100000", x"ae8d0000", x"85644e78", x"c2f6b9b0", x"a78a1f4c", x"c7ef3d40"),
	(x"fd7201b5", x"4ff70000", x"24a60000", x"7a930000", x"70060dad", x"6d27dc98", x"975a4af4", x"f78c5d47", x"1aa30188", x"5feb8000", x"98ec0000", x"38560000", x"bfef2385", x"293c1743", x"8be758c3", x"6b6151c8"),
	(x"ad8d01b1", x"0a834000", x"195d0000", x"63750000", x"6bba5bab", x"8c55a7c5", x"76f28662", x"8c978bfe", x"ec23018d", x"6ba84000", x"bceb0000", x"b76b0000", x"9ed8187e", x"2384c2ed", x"4622d3da", x"bcf4ebf9"),
	(x"5b0d01b4", x"3ec08000", x"3d5a0000", x"ec480000", x"4a8d6050", x"86ed726b", x"bb370d7b", x"5b0231cf", x"4a5c018c", x"1a9fc000", x"a5170000", x"21b00000", x"a4537583", x"c84e6c1e", x"6a4f9455", x"107a8771"),
	(x"fc8701b9", x"b4880000", x"c3770000", x"f13c0000", x"53a42fff", x"9f773f8c", x"201830a3", x"be0f7f6c", x"68b60189", x"a314c000", x"24bf0000", x"e4a40000", x"792a0c02", x"0b423fdc", x"3fbc8948", x"30a9fe60"),
	(x"0a0701bc", x"80cbc000", x"e7700000", x"7e010000", x"72931404", x"95cfea22", x"edddbbba", x"699ac55d", x"cec90188", x"d2234000", x"3d430000", x"727f0000", x"43a161ff", x"e088912f", x"13d1cec7", x"9c2792e8"),
	(x"5af801b8", x"c5bf8000", x"da8b0000", x"67e70000", x"692f4202", x"74bd917f", x"0c75772c", x"128113e4", x"3849018d", x"e6608000", x"19440000", x"fd420000", x"62965a04", x"ea304481", x"de1445de", x"4bb228d9"),
	(x"ac7801bd", x"f1fc4000", x"fe8c0000", x"e8da0000", x"481879f9", x"7e0544d1", x"c1b0fc35", x"c514a9d5", x"9e36018c", x"97570000", x"00b80000", x"6b990000", x"581d37f9", x"01faea72", x"f2790251", x"e73c4451")
    ),(
	(x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000"),
	(x"0c720000", x"49e50f00", x"42790000", x"5cea0000", x"33aa301a", x"15822514", x"95a34b7b", x"b44b0090", x"fe220000", x"a7580500", x"25d10000", x"f7600000", x"893178da", x"1fd4f860", x"4ed0a315", x"a123ff9f"),
	(x"fe220000", x"a7580500", x"25d10000", x"f7600000", x"893178da", x"1fd4f860", x"4ed0a315", x"a123ff9f", x"f2500000", x"eebd0a00", x"67a80000", x"ab8a0000", x"ba9b48c0", x"0a56dd74", x"db73e86e", x"1568ff0f"),
	(x"f2500000", x"eebd0a00", x"67a80000", x"ab8a0000", x"ba9b48c0", x"0a56dd74", x"db73e86e", x"1568ff0f", x"0c720000", x"49e50f00", x"42790000", x"5cea0000", x"33aa301a", x"15822514", x"95a34b7b", x"b44b0090"),
	(x"45180000", x"a5b51700", x"f96a0000", x"3b480000", x"1ecc142c", x"231395d6", x"16bca6b0", x"df33f4df", x"b83d0000", x"16710600", x"379a0000", x"f5b10000", x"228161ac", x"ae48f145", x"66241616", x"c5c1eb3e"),
	(x"496a0000", x"ec501800", x"bb130000", x"67a20000", x"2d662436", x"3691b0c2", x"831fedcb", x"6b78f44f", x"461f0000", x"b1290300", x"124b0000", x"02d10000", x"abb01976", x"b19c0925", x"28f4b503", x"64e214a1"),
	(x"bb3a0000", x"02ed1200", x"dcbb0000", x"cc280000", x"97fd6cf6", x"3cc76db6", x"586c05a5", x"7e100b40", x"4a6d0000", x"f8cc0c00", x"50320000", x"5e3b0000", x"981a296c", x"a41e2c31", x"bd57fe78", x"d0a91431"),
	(x"b7480000", x"4b081d00", x"9ec20000", x"90c20000", x"a4575cec", x"294548a2", x"cdcf4ede", x"ca5b0bd0", x"b44f0000", x"5f940900", x"75e30000", x"a95b0000", x"112b51b6", x"bbcad451", x"f3875d6d", x"718aebae"),
	(x"b83d0000", x"16710600", x"379a0000", x"f5b10000", x"228161ac", x"ae48f145", x"66241616", x"c5c1eb3e", x"fd250000", x"b3c41100", x"cef00000", x"cef90000", x"3c4d7580", x"8d5b6493", x"7098b0a6", x"1af21fe1"),
	(x"b44f0000", x"5f940900", x"75e30000", x"a95b0000", x"112b51b6", x"bbcad451", x"f3875d6d", x"718aebae", x"03070000", x"149c1400", x"eb210000", x"39990000", x"b57c0d5a", x"928f9cf3", x"3e4813b3", x"bbd1e07e"),
	(x"461f0000", x"b1290300", x"124b0000", x"02d10000", x"abb01976", x"b19c0925", x"28f4b503", x"64e214a1", x"0f750000", x"5d791b00", x"a9580000", x"65730000", x"86d63d40", x"870db9e7", x"abeb58c8", x"0f9ae0ee"),
	(x"4a6d0000", x"f8cc0c00", x"50320000", x"5e3b0000", x"981a296c", x"a41e2c31", x"bd57fe78", x"d0a91431", x"f1570000", x"fa211e00", x"8c890000", x"92130000", x"0fe7459a", x"98d94187", x"e53bfbdd", x"aeb91f71"),
	(x"fd250000", x"b3c41100", x"cef00000", x"cef90000", x"3c4d7580", x"8d5b6493", x"7098b0a6", x"1af21fe1", x"45180000", x"a5b51700", x"f96a0000", x"3b480000", x"1ecc142c", x"231395d6", x"16bca6b0", x"df33f4df"),
	(x"f1570000", x"fa211e00", x"8c890000", x"92130000", x"0fe7459a", x"98d94187", x"e53bfbdd", x"aeb91f71", x"bb3a0000", x"02ed1200", x"dcbb0000", x"cc280000", x"97fd6cf6", x"3cc76db6", x"586c05a5", x"7e100b40"),
	(x"03070000", x"149c1400", x"eb210000", x"39990000", x"b57c0d5a", x"928f9cf3", x"3e4813b3", x"bbd1e07e", x"b7480000", x"4b081d00", x"9ec20000", x"90c20000", x"a4575cec", x"294548a2", x"cdcf4ede", x"ca5b0bd0"),
	(x"0f750000", x"5d791b00", x"a9580000", x"65730000", x"86d63d40", x"870db9e7", x"abeb58c8", x"0f9ae0ee", x"496a0000", x"ec501800", x"bb130000", x"67a20000", x"2d662436", x"3691b0c2", x"831fedcb", x"6b78f44f"),
	(x"75a40000", x"c28b2700", x"94a40000", x"90f50000", x"fb7857e0", x"49ce0bae", x"1767c483", x"aedf667e", x"d1660000", x"1bbc0300", x"9eec0000", x"f6940000", x"03024527", x"cf70fcf2", x"b4431b17", x"857f3c2b"),
	(x"79d60000", x"8b6e2800", x"d6dd0000", x"cc1f0000", x"c8d267fa", x"5c4c2eba", x"82c48ff8", x"1a9466ee", x"2f440000", x"bce40600", x"bb3d0000", x"01f40000", x"8a333dfd", x"d0a40492", x"fa93b802", x"245cc3b4"),
	(x"8b860000", x"65d32200", x"b1750000", x"67950000", x"72492f3a", x"561af3ce", x"59b76796", x"0ffc99e1", x"23360000", x"f5010900", x"f9440000", x"5d1e0000", x"b9990de7", x"c5262186", x"6f30f379", x"9017c324"),
	(x"87f40000", x"2c362d00", x"f30c0000", x"3b7f0000", x"41e31f20", x"4398d6da", x"cc142ced", x"bbb79971", x"dd140000", x"52590c00", x"dc950000", x"aa7e0000", x"30a8753d", x"daf2d9e6", x"21e0506c", x"31343cbb"),
	(x"30bc0000", x"673e3000", x"6dce0000", x"abbd0000", x"e5b443cc", x"6add9e78", x"01db6233", x"71ec92a1", x"695b0000", x"0dcd0500", x"a9760000", x"03250000", x"2183248b", x"61380db7", x"d2670d01", x"40bed715"),
	(x"3cce0000", x"2edb3f00", x"2fb70000", x"f7570000", x"d61e73d6", x"7f5fbb6c", x"94782948", x"c5a79231", x"97790000", x"aa950000", x"8ca70000", x"f4450000", x"a8b25c51", x"7eecf5d7", x"9cb7ae14", x"e19d288a"),
	(x"ce9e0000", x"c0663500", x"481f0000", x"5cdd0000", x"6c853b16", x"75096618", x"4f0bc126", x"d0cf6d3e", x"9b0b0000", x"e3700f00", x"cede0000", x"a8af0000", x"9b186c4b", x"6b6ed0c3", x"0914e56f", x"55d6281a"),
	(x"c2ec0000", x"89833a00", x"0a660000", x"00370000", x"5f2f0b0c", x"608b430c", x"daa88a5d", x"64846dae", x"65290000", x"44280a00", x"eb0f0000", x"5fcf0000", x"12291491", x"74ba28a3", x"47c4467a", x"f4f5d785"),
	(x"cd990000", x"d4fa2100", x"a33e0000", x"65440000", x"d9f9364c", x"e786faeb", x"7143d295", x"6b1e8d40", x"2c430000", x"a8781200", x"501c0000", x"386d0000", x"3f4f30a7", x"422b9861", x"c4dbabb1", x"9f8d23ca"),
	(x"c1eb0000", x"9d1f2e00", x"e1470000", x"39ae0000", x"ea530656", x"f204dfff", x"e4e099ee", x"df558dd0", x"d2610000", x"0f201700", x"75cd0000", x"cf0d0000", x"b67e487d", x"5dff6001", x"8a0b08a4", x"3eaedc55"),
	(x"33bb0000", x"73a22400", x"86ef0000", x"92240000", x"50c84e96", x"f852028b", x"3f937180", x"ca3d72df", x"de130000", x"46c51800", x"37b40000", x"93e70000", x"85d47867", x"487d4515", x"1fa843df", x"8ae5dcc5"),
	(x"3fc90000", x"3a472b00", x"c4960000", x"cece0000", x"63627e8c", x"edd0279f", x"aa303afb", x"7e76724f", x"20310000", x"e19d1d00", x"12650000", x"64870000", x"0ce500bd", x"57a9bd75", x"5178e0ca", x"2bc6235a"),
	(x"88810000", x"714f3600", x"5a540000", x"5e0c0000", x"c7352260", x"c4956f3d", x"67ff7425", x"b42d799f", x"947e0000", x"be091400", x"67860000", x"cddc0000", x"1dce510b", x"ec636924", x"a2ffbda7", x"5a4cc8f4"),
	(x"84f30000", x"38aa3900", x"182d0000", x"02e60000", x"f49f127a", x"d1174a29", x"f25c3f5e", x"0066790f", x"6a5c0000", x"19511100", x"42570000", x"3abc0000", x"94ff29d1", x"f3b79144", x"ec2f1eb2", x"fb6f376b"),
	(x"76a30000", x"d6173300", x"7f850000", x"a96c0000", x"4e045aba", x"db41975d", x"292fd730", x"150e8600", x"662e0000", x"50b41e00", x"002e0000", x"66560000", x"a75519cb", x"e635b450", x"798c55c9", x"4f2437fb"),
	(x"7ad10000", x"9ff23c00", x"3dfc0000", x"f5860000", x"7dae6aa0", x"cec3b249", x"bc8c9c4b", x"a1458690", x"980c0000", x"f7ec1b00", x"25ff0000", x"91360000", x"2e646111", x"f9e14c30", x"375cf6dc", x"ee07c864"),
	(x"d1660000", x"1bbc0300", x"9eec0000", x"f6940000", x"03024527", x"cf70fcf2", x"b4431b17", x"857f3c2b", x"a4c20000", x"d9372400", x"0a480000", x"66610000", x"f87a12c7", x"86bef75c", x"a324df94", x"2ba05a55"),
	(x"dd140000", x"52590c00", x"dc950000", x"aa7e0000", x"30a8753d", x"daf2d9e6", x"21e0506c", x"31343cbb", x"5ae00000", x"7e6f2100", x"2f990000", x"91010000", x"714b6a1d", x"996a0f3c", x"edf47c81", x"8a83a5ca"),
	(x"2f440000", x"bce40600", x"bb3d0000", x"01f40000", x"8a333dfd", x"d0a40492", x"fa93b802", x"245cc3b4", x"56920000", x"378a2e00", x"6de00000", x"cdeb0000", x"42e15a07", x"8ce82a28", x"785737fa", x"3ec8a55a"),
	(x"23360000", x"f5010900", x"f9440000", x"5d1e0000", x"b9990de7", x"c5262186", x"6f30f379", x"9017c324", x"a8b00000", x"90d22b00", x"48310000", x"3a8b0000", x"cbd022dd", x"933cd248", x"368794ef", x"9feb5ac5"),
	(x"947e0000", x"be091400", x"67860000", x"cddc0000", x"1dce510b", x"ec636924", x"a2ffbda7", x"5a4cc8f4", x"1cff0000", x"cf462200", x"3dd20000", x"93d00000", x"dafb736b", x"28f60619", x"c500c982", x"ee61b16b"),
	(x"980c0000", x"f7ec1b00", x"25ff0000", x"91360000", x"2e646111", x"f9e14c30", x"375cf6dc", x"ee07c864", x"e2dd0000", x"681e2700", x"18030000", x"64b00000", x"53ca0bb1", x"3722fe79", x"8bd06a97", x"4f424ef4"),
	(x"6a5c0000", x"19511100", x"42570000", x"3abc0000", x"94ff29d1", x"f3b79144", x"ec2f1eb2", x"fb6f376b", x"eeaf0000", x"21fb2800", x"5a7a0000", x"385a0000", x"60603bab", x"22a0db6d", x"1e7321ec", x"fb094e64"),
	(x"662e0000", x"50b41e00", x"002e0000", x"66560000", x"a75519cb", x"e635b450", x"798c55c9", x"4f2437fb", x"108d0000", x"86a32d00", x"7fab0000", x"cf3a0000", x"e9514371", x"3d74230d", x"50a382f9", x"5a2ab1fb"),
	(x"695b0000", x"0dcd0500", x"a9760000", x"03250000", x"2183248b", x"61380db7", x"d2670d01", x"40bed715", x"59e70000", x"6af33500", x"c4b80000", x"a8980000", x"c4376747", x"0be593cf", x"d3bc6f32", x"315245b4"),
	(x"65290000", x"44280a00", x"eb0f0000", x"5fcf0000", x"12291491", x"74ba28a3", x"47c4467a", x"f4f5d785", x"a7c50000", x"cdab3000", x"e1690000", x"5ff80000", x"4d061f9d", x"14316baf", x"9d6ccc27", x"9071ba2b"),
	(x"97790000", x"aa950000", x"8ca70000", x"f4450000", x"a8b25c51", x"7eecf5d7", x"9cb7ae14", x"e19d288a", x"abb70000", x"844e3f00", x"a3100000", x"03120000", x"7eac2f87", x"01b34ebb", x"08cf875c", x"243ababb"),
	(x"9b0b0000", x"e3700f00", x"cede0000", x"a8af0000", x"9b186c4b", x"6b6ed0c3", x"0914e56f", x"55d6281a", x"55950000", x"23163a00", x"86c10000", x"f4720000", x"f79d575d", x"1e67b6db", x"461f2449", x"85194524"),
	(x"2c430000", x"a8781200", x"501c0000", x"386d0000", x"3f4f30a7", x"422b9861", x"c4dbabb1", x"9f8d23ca", x"e1da0000", x"7c823300", x"f3220000", x"5d290000", x"e6b606eb", x"a5ad628a", x"b5987924", x"f493ae8a"),
	(x"20310000", x"e19d1d00", x"12650000", x"64870000", x"0ce500bd", x"57a9bd75", x"5178e0ca", x"2bc6235a", x"1ff80000", x"dbda3600", x"d6f30000", x"aa490000", x"6f877e31", x"ba799aea", x"fb48da31", x"55b05115"),
	(x"d2610000", x"0f201700", x"75cd0000", x"cf0d0000", x"b67e487d", x"5dff6001", x"8a0b08a4", x"3eaedc55", x"138a0000", x"923f3900", x"948a0000", x"f6a30000", x"5c2d4e2b", x"affbbffe", x"6eeb914a", x"e1fb5185"),
	(x"de130000", x"46c51800", x"37b40000", x"93e70000", x"85d47867", x"487d4515", x"1fa843df", x"8ae5dcc5", x"eda80000", x"35673c00", x"b15b0000", x"01c30000", x"d51c36f1", x"b02f479e", x"203b325f", x"40d8ae1a"),
	(x"a4c20000", x"d9372400", x"0a480000", x"66610000", x"f87a12c7", x"86bef75c", x"a324df94", x"2ba05a55", x"75a40000", x"c28b2700", x"94a40000", x"90f50000", x"fb7857e0", x"49ce0bae", x"1767c483", x"aedf667e"),
	(x"a8b00000", x"90d22b00", x"48310000", x"3a8b0000", x"cbd022dd", x"933cd248", x"368794ef", x"9feb5ac5", x"8b860000", x"65d32200", x"b1750000", x"67950000", x"72492f3a", x"561af3ce", x"59b76796", x"0ffc99e1"),
	(x"5ae00000", x"7e6f2100", x"2f990000", x"91010000", x"714b6a1d", x"996a0f3c", x"edf47c81", x"8a83a5ca", x"87f40000", x"2c362d00", x"f30c0000", x"3b7f0000", x"41e31f20", x"4398d6da", x"cc142ced", x"bbb79971"),
	(x"56920000", x"378a2e00", x"6de00000", x"cdeb0000", x"42e15a07", x"8ce82a28", x"785737fa", x"3ec8a55a", x"79d60000", x"8b6e2800", x"d6dd0000", x"cc1f0000", x"c8d267fa", x"5c4c2eba", x"82c48ff8", x"1a9466ee"),
	(x"e1da0000", x"7c823300", x"f3220000", x"5d290000", x"e6b606eb", x"a5ad628a", x"b5987924", x"f493ae8a", x"cd990000", x"d4fa2100", x"a33e0000", x"65440000", x"d9f9364c", x"e786faeb", x"7143d295", x"6b1e8d40"),
	(x"eda80000", x"35673c00", x"b15b0000", x"01c30000", x"d51c36f1", x"b02f479e", x"203b325f", x"40d8ae1a", x"33bb0000", x"73a22400", x"86ef0000", x"92240000", x"50c84e96", x"f852028b", x"3f937180", x"ca3d72df"),
	(x"1ff80000", x"dbda3600", x"d6f30000", x"aa490000", x"6f877e31", x"ba799aea", x"fb48da31", x"55b05115", x"3fc90000", x"3a472b00", x"c4960000", x"cece0000", x"63627e8c", x"edd0279f", x"aa303afb", x"7e76724f"),
	(x"138a0000", x"923f3900", x"948a0000", x"f6a30000", x"5c2d4e2b", x"affbbffe", x"6eeb914a", x"e1fb5185", x"c1eb0000", x"9d1f2e00", x"e1470000", x"39ae0000", x"ea530656", x"f204dfff", x"e4e099ee", x"df558dd0"),
	(x"1cff0000", x"cf462200", x"3dd20000", x"93d00000", x"dafb736b", x"28f60619", x"c500c982", x"ee61b16b", x"88810000", x"714f3600", x"5a540000", x"5e0c0000", x"c7352260", x"c4956f3d", x"67ff7425", x"b42d799f"),
	(x"108d0000", x"86a32d00", x"7fab0000", x"cf3a0000", x"e9514371", x"3d74230d", x"50a382f9", x"5a2ab1fb", x"76a30000", x"d6173300", x"7f850000", x"a96c0000", x"4e045aba", x"db41975d", x"292fd730", x"150e8600"),
	(x"e2dd0000", x"681e2700", x"18030000", x"64b00000", x"53ca0bb1", x"3722fe79", x"8bd06a97", x"4f424ef4", x"7ad10000", x"9ff23c00", x"3dfc0000", x"f5860000", x"7dae6aa0", x"cec3b249", x"bc8c9c4b", x"a1458690"),
	(x"eeaf0000", x"21fb2800", x"5a7a0000", x"385a0000", x"60603bab", x"22a0db6d", x"1e7321ec", x"fb094e64", x"84f30000", x"38aa3900", x"182d0000", x"02e60000", x"f49f127a", x"d1174a29", x"f25c3f5e", x"0066790f"),
	(x"59e70000", x"6af33500", x"c4b80000", x"a8980000", x"c4376747", x"0be593cf", x"d3bc6f32", x"315245b4", x"30bc0000", x"673e3000", x"6dce0000", x"abbd0000", x"e5b443cc", x"6add9e78", x"01db6233", x"71ec92a1"),
	(x"55950000", x"23163a00", x"86c10000", x"f4720000", x"f79d575d", x"1e67b6db", x"461f2449", x"85194524", x"ce9e0000", x"c0663500", x"481f0000", x"5cdd0000", x"6c853b16", x"75096618", x"4f0bc126", x"d0cf6d3e"),
	(x"a7c50000", x"cdab3000", x"e1690000", x"5ff80000", x"4d061f9d", x"14316baf", x"9d6ccc27", x"9071ba2b", x"c2ec0000", x"89833a00", x"0a660000", x"00370000", x"5f2f0b0c", x"608b430c", x"daa88a5d", x"64846dae"),
	(x"abb70000", x"844e3f00", x"a3100000", x"03120000", x"7eac2f87", x"01b34ebb", x"08cf875c", x"243ababb", x"3cce0000", x"2edb3f00", x"2fb70000", x"f7570000", x"d61e73d6", x"7f5fbb6c", x"94782948", x"c5a79231"),
	(x"75c90003", x"0e10c000", x"d1200000", x"baea0000", x"8bc42f3e", x"8758b757", x"bb28761d", x"00b72e2b", x"eecf0001", x"6f564000", x"f33e0000", x"a79e0000", x"bdb57219", x"b711ebc5", x"4a3b40ba", x"feabf254"),
	(x"79bb0003", x"47f5cf00", x"93590000", x"e6000000", x"b86e1f24", x"92da9243", x"2e8b3d66", x"b4fc2ebb", x"10ed0001", x"c80e4500", x"d6ef0000", x"50fe0000", x"34840ac3", x"a8c513a5", x"04ebe3af", x"5f880dcb"),
	(x"8beb0003", x"a948c500", x"f4f10000", x"4d8a0000", x"02f557e4", x"988c4f37", x"f5f8d508", x"a194d1b4", x"1c9f0001", x"81eb4a00", x"94960000", x"0c140000", x"072e3ad9", x"bd4736b1", x"9148a8d4", x"ebc30d5b"),
	(x"87990003", x"e0adca00", x"b6880000", x"11600000", x"315f67fe", x"8d0e6a23", x"605b9e73", x"15dfd124", x"e2bd0001", x"26b34f00", x"b1470000", x"fb740000", x"8e1f4203", x"a293ced1", x"df980bc1", x"4ae0f2c4"),
	(x"30d10003", x"aba5d700", x"284a0000", x"81a20000", x"95083b12", x"a44b2281", x"ad94d0ad", x"df84daf4", x"56f20001", x"79274600", x"c4a40000", x"522f0000", x"9f3413b5", x"19591a80", x"2c1f56ac", x"3b6a196a"),
	(x"3ca30003", x"e240d800", x"6a330000", x"dd480000", x"a6a20b08", x"b1c90795", x"38379bd6", x"6bcfda64", x"a8d00001", x"de7f4300", x"e1750000", x"a54f0000", x"16056b6f", x"068de2e0", x"62cff5b9", x"9a49e6f5"),
	(x"cef30003", x"0cfdd200", x"0d9b0000", x"76c20000", x"1c3943c8", x"bb9fdae1", x"e34473b8", x"7ea7256b", x"a4a20001", x"979a4c00", x"a30c0000", x"f9a50000", x"25af5b75", x"130fc7f4", x"f76cbec2", x"2e02e665"),
	(x"c2810003", x"4518dd00", x"4fe20000", x"2a280000", x"2f9373d2", x"ae1dfff5", x"76e738c3", x"caec25fb", x"5a800001", x"30c24900", x"86dd0000", x"0ec50000", x"ac9e23af", x"0cdb3f94", x"b9bc1dd7", x"8f2119fa"),
	(x"cdf40003", x"1861c600", x"e6ba0000", x"4f5b0000", x"a9454e92", x"29104612", x"dd0c600b", x"c576c515", x"13ea0001", x"dc925100", x"3dce0000", x"69670000", x"81f80799", x"3a4a8f56", x"3aa3f01c", x"e459edb5"),
	(x"c1860003", x"5184c900", x"a4c30000", x"13b10000", x"9aef7e88", x"3c926306", x"48af2b70", x"713dc585", x"edc80001", x"7bca5400", x"181f0000", x"9e070000", x"08c97f43", x"259e7736", x"74735309", x"457a122a"),
	(x"33d60003", x"bf39c300", x"c36b0000", x"b83b0000", x"20743648", x"36c4be72", x"93dcc31e", x"64553a8a", x"e1ba0001", x"322f5b00", x"5a660000", x"c2ed0000", x"3b634f59", x"301c5222", x"e1d01872", x"f13112ba"),
	(x"3fa40003", x"f6dccc00", x"81120000", x"e4d10000", x"13de0652", x"23469b66", x"067f8865", x"d01e3a1a", x"1f980001", x"95775e00", x"7fb70000", x"358d0000", x"b2523783", x"2fc8aa42", x"af00bb67", x"5012ed25"),
	(x"88ec0003", x"bdd4d100", x"1fd00000", x"74130000", x"b7895abe", x"0a03d3c4", x"cbb0c6bb", x"1a4531ca", x"abd70001", x"cae35700", x"0a540000", x"9cd60000", x"a3796635", x"94027e13", x"5c87e60a", x"2198068b"),
	(x"849e0003", x"f431de00", x"5da90000", x"28f90000", x"84236aa4", x"1f81f6d0", x"5e138dc0", x"ae0e315a", x"55f50001", x"6dbb5200", x"2f850000", x"6bb60000", x"2a481eef", x"8bd68673", x"1257451f", x"80bbf914"),
	(x"76ce0003", x"1a8cd400", x"3a010000", x"83730000", x"3eb82264", x"15d72ba4", x"856065ae", x"bb66ce55", x"59870001", x"245e5d00", x"6dfc0000", x"375c0000", x"19e22ef5", x"9e54a367", x"87f40e64", x"34f0f984"),
	(x"7abc0003", x"5369db00", x"78780000", x"df990000", x"0d12127e", x"00550eb0", x"10c32ed5", x"0f2dcec5", x"a7a50001", x"83065800", x"482d0000", x"c03c0000", x"90d3562f", x"81805b07", x"c924ad71", x"95d3061b"),
	(x"006d0003", x"cc9be700", x"45840000", x"2a1f0000", x"70bc78de", x"ce96bcf9", x"ac4fb29e", x"ae684855", x"3fa90001", x"74ea4300", x"6dd20000", x"510a0000", x"beb7373e", x"78611737", x"fe785bad", x"7bd4ce7f"),
	(x"0c1f0003", x"857ee800", x"07fd0000", x"76f50000", x"431648c4", x"db1499ed", x"39ecf9e5", x"1a2348c5", x"c18b0001", x"d3b24600", x"48030000", x"a66a0000", x"37864fe4", x"67b5ef57", x"b0a8f8b8", x"daf731e0"),
	(x"fe4f0003", x"6bc3e200", x"60550000", x"dd7f0000", x"f98d0004", x"d1424499", x"e29f118b", x"0f4bb7ca", x"cdf90001", x"9a574900", x"0a7a0000", x"fa800000", x"042c7ffe", x"7237ca43", x"250bb3c3", x"6ebc3170"),
	(x"f23d0003", x"2226ed00", x"222c0000", x"81950000", x"ca27301e", x"c4c0618d", x"773c5af0", x"bb00b75a", x"33db0001", x"3d0f4c00", x"2fab0000", x"0de00000", x"8d1d0724", x"6de33223", x"6bdb10d6", x"cf9fceef"),
	(x"45750003", x"692ef000", x"bcee0000", x"11570000", x"6e706cf2", x"ed85292f", x"baf3142e", x"715bbc8a", x"87940001", x"629b4500", x"5a480000", x"a4bb0000", x"9c365692", x"d629e672", x"985c4dbb", x"be152541"),
	(x"49070003", x"20cbff00", x"fe970000", x"4dbd0000", x"5dda5ce8", x"f8070c3b", x"2f505f55", x"c510bc1a", x"79b60001", x"c5c34000", x"7f990000", x"53db0000", x"15072e48", x"c9fd1e12", x"d68ceeae", x"1f36dade"),
	(x"bb570003", x"ce76f500", x"993f0000", x"e6370000", x"e7411428", x"f251d14f", x"f423b73b", x"d0784315", x"75c40001", x"8c264f00", x"3de00000", x"0f310000", x"26ad1e52", x"dc7f3b06", x"432fa5d5", x"ab7dda4e"),
	(x"b7250003", x"8793fa00", x"db460000", x"badd0000", x"d4eb2432", x"e7d3f45b", x"6180fc40", x"64334385", x"8be60001", x"2b7e4a00", x"18310000", x"f8510000", x"af9c6688", x"c3abc366", x"0dff06c0", x"0a5e25d1"),
	(x"b8500003", x"daeae100", x"721e0000", x"dfae0000", x"523d1972", x"60de4dbc", x"ca6ba488", x"6ba9a36b", x"c28c0001", x"c72e5200", x"a3220000", x"9ff30000", x"82fa42be", x"f53a73a4", x"8ee0eb0b", x"6126d19e"),
	(x"b4220003", x"930fee00", x"30670000", x"83440000", x"61972968", x"755c68a8", x"5fc8eff3", x"dfe2a3fb", x"3cae0001", x"60765700", x"86f30000", x"68930000", x"0bcb3a64", x"eaee8bc4", x"c030481e", x"c0052e01"),
	(x"46720003", x"7db2e400", x"57cf0000", x"28ce0000", x"db0c61a8", x"7f0ab5dc", x"84bb079d", x"ca8a5cf4", x"30dc0001", x"29935800", x"c48a0000", x"34790000", x"38610a7e", x"ff6caed0", x"55930365", x"744e2e91"),
	(x"4a000003", x"3457eb00", x"15b60000", x"74240000", x"e8a651b2", x"6a8890c8", x"11184ce6", x"7ec15c64", x"cefe0001", x"8ecb5d00", x"e15b0000", x"c3190000", x"b15072a4", x"e0b856b0", x"1b43a070", x"d56dd10e"),
	(x"fd480003", x"7f5ff600", x"8b740000", x"e4e60000", x"4cf10d5e", x"43cdd86a", x"dcd70238", x"b49a57b4", x"7ab10001", x"d15f5400", x"94b80000", x"6a420000", x"a07b2312", x"5b7282e1", x"e8c4fd1d", x"a4e73aa0"),
	(x"f13a0003", x"36baf900", x"c90d0000", x"b80c0000", x"7f5b3d44", x"564ffd7e", x"49744943", x"00d15724", x"84930001", x"76075100", x"b1690000", x"9d220000", x"294a5bc8", x"44a67a81", x"a6145e08", x"05c4c53f"),
	(x"036a0003", x"d807f300", x"aea50000", x"13860000", x"c5c07584", x"5c19200a", x"9207a12d", x"15b9a82b", x"88e10001", x"3fe25e00", x"f3100000", x"c1c80000", x"1ae06bd2", x"51245f95", x"33b71573", x"b18fc5af"),
	(x"0f180003", x"91e2fc00", x"ecdc0000", x"4f6c0000", x"f66a459e", x"499b051e", x"07a4ea56", x"a1f2a8bb", x"76c30001", x"98ba5b00", x"d6c10000", x"36a80000", x"93d11308", x"4ef0a7f5", x"7d67b666", x"10ac3a30"),
	(x"a4af0003", x"15acc300", x"4fcc0000", x"4c7e0000", x"88c66a19", x"48284ba5", x"0f6b6d0a", x"85c81200", x"4a0d0001", x"b6616400", x"f9760000", x"c1ff0000", x"45cf60de", x"31af1c99", x"e91f9f2e", x"d50ba801"),
	(x"a8dd0003", x"5c49cc00", x"0db50000", x"10940000", x"bb6c5a03", x"5daa6eb1", x"9ac82671", x"31831290", x"b42f0001", x"11396100", x"dca70000", x"369f0000", x"ccfe1804", x"2e7be4f9", x"a7cf3c3b", x"7428579e"),
	(x"5a8d0003", x"b2f4c600", x"6a1d0000", x"bb1e0000", x"01f712c3", x"57fcb3c5", x"41bbce1f", x"24ebed9f", x"b85d0001", x"58dc6e00", x"9ede0000", x"6a750000", x"ff54281e", x"3bf9c1ed", x"326c7740", x"c063570e"),
	(x"56ff0003", x"fb11c900", x"28640000", x"e7f40000", x"325d22d9", x"427e96d1", x"d4188564", x"90a0ed0f", x"467f0001", x"ff846b00", x"bb0f0000", x"9d150000", x"766550c4", x"242d398d", x"7cbcd455", x"6140a891"),
	(x"e1b70003", x"b019d400", x"b6a60000", x"77360000", x"960a7e35", x"6b3bde73", x"19d7cbba", x"5afbe6df", x"f2300001", x"a0106200", x"ceec0000", x"344e0000", x"674e0172", x"9fe7eddc", x"8f3b8938", x"10ca433f"),
	(x"edc50003", x"f9fcdb00", x"f4df0000", x"2bdc0000", x"a5a04e2f", x"7eb9fb67", x"8c7480c1", x"eeb0e64f", x"0c120001", x"07486700", x"eb3d0000", x"c32e0000", x"ee7f79a8", x"803315bc", x"c1eb2a2d", x"b1e9bca0"),
	(x"1f950003", x"1741d100", x"93770000", x"80560000", x"1f3b06ef", x"74ef2613", x"570768af", x"fbd81940", x"00600001", x"4ead6800", x"a9440000", x"9fc40000", x"ddd549b2", x"95b130a8", x"54486156", x"05a2bc30"),
	(x"13e70003", x"5ea4de00", x"d10e0000", x"dcbc0000", x"2c9136f5", x"616d0307", x"c2a423d4", x"4f9319d0", x"fe420001", x"e9f56d00", x"8c950000", x"68a40000", x"54e43168", x"8a65c8c8", x"1a98c243", x"a48143af"),
	(x"1c920003", x"03ddc500", x"78560000", x"b9cf0000", x"aa470bb5", x"e660bae0", x"694f7b1c", x"4009f93e", x"b7280001", x"05a57500", x"37860000", x"0f060000", x"7982155e", x"bcf4780a", x"99872f88", x"cff9b7e0"),
	(x"10e00003", x"4a38ca00", x"3a2f0000", x"e5250000", x"99ed3baf", x"f3e29ff4", x"fcec3067", x"f442f9ae", x"490a0001", x"a2fd7000", x"12570000", x"f8660000", x"f0b36d84", x"a320806a", x"d7578c9d", x"6eda487f"),
	(x"e2b00003", x"a485c000", x"5d870000", x"4eaf0000", x"2376736f", x"f9b44280", x"279fd809", x"e12a06a1", x"45780001", x"eb187f00", x"502e0000", x"a48c0000", x"c3195d9e", x"b6a2a57e", x"42f4c7e6", x"da9148ef"),
	(x"eec20003", x"ed60cf00", x"1ffe0000", x"12450000", x"10dc4375", x"ec366794", x"b23c9372", x"55610631", x"bb5a0001", x"4c407a00", x"75ff0000", x"53ec0000", x"4a282544", x"a9765d1e", x"0c2464f3", x"7bb2b770"),
	(x"598a0003", x"a668d200", x"813c0000", x"82870000", x"b48b1f99", x"c5732f36", x"7ff3ddac", x"9f3a0de1", x"0f150001", x"13d47300", x"001c0000", x"fab70000", x"5b0374f2", x"12bc894f", x"ffa3399e", x"0a385cde"),
	(x"55f80003", x"ef8ddd00", x"c3450000", x"de6d0000", x"87212f83", x"d0f10a22", x"ea5096d7", x"2b710d71", x"f1370001", x"b48c7600", x"25cd0000", x"0dd70000", x"d2320c28", x"0d68712f", x"b1739a8b", x"ab1ba341"),
	(x"a7a80003", x"0130d700", x"a4ed0000", x"75e70000", x"3dba6743", x"daa7d756", x"31237eb9", x"3e19f27e", x"fd450001", x"fd697900", x"67b40000", x"513d0000", x"e1983c32", x"18ea543b", x"24d0d1f0", x"1f50a3d1"),
	(x"abda0003", x"48d5d800", x"e6940000", x"290d0000", x"0e105759", x"cf25f242", x"a48035c2", x"8a52f2ee", x"03670001", x"5a317c00", x"42650000", x"a65d0000", x"68a944e8", x"073eac5b", x"6a0072e5", x"be735c4e"),
	(x"d10b0003", x"d727e400", x"db680000", x"dc8b0000", x"73be3df9", x"01e6400b", x"180ca989", x"2b17747e", x"9b6b0001", x"addd6700", x"679a0000", x"376b0000", x"46cd25f9", x"fedfe06b", x"5d5c8439", x"5074942a"),
	(x"dd790003", x"9ec2eb00", x"99110000", x"80610000", x"40140de3", x"1464651f", x"8dafe2f2", x"9f5c74ee", x"65490001", x"0a856200", x"424b0000", x"c00b0000", x"cffc5d23", x"e10b180b", x"138c272c", x"f1576bb5"),
	(x"2f290003", x"707fe100", x"feb90000", x"2beb0000", x"fa8f4523", x"1e32b86b", x"56dc0a9c", x"8a348be1", x"693b0001", x"43606d00", x"00320000", x"9ce10000", x"fc566d39", x"f4893d1f", x"862f6c57", x"451c6b25"),
	(x"235b0003", x"399aee00", x"bcc00000", x"77010000", x"c9257539", x"0bb09d7f", x"c37f41e7", x"3e7f8b71", x"97190001", x"e4386800", x"25e30000", x"6b810000", x"756715e3", x"eb5dc57f", x"c8ffcf42", x"e43f94ba"),
	(x"94130003", x"7292f300", x"22020000", x"e7c30000", x"6d7229d5", x"22f5d5dd", x"0eb00f39", x"f42480a1", x"23560001", x"bbac6100", x"50000000", x"c2da0000", x"644c4455", x"5097112e", x"3b78922f", x"95b57f14"),
	(x"98610003", x"3b77fc00", x"607b0000", x"bb290000", x"5ed819cf", x"3777f0c9", x"9b134442", x"406f8031", x"dd740001", x"1cf46400", x"75d10000", x"35ba0000", x"ed7d3c8f", x"4f43e94e", x"75a8313a", x"3496808b"),
	(x"6a310003", x"d5caf600", x"07d30000", x"10a30000", x"e443510f", x"3d212dbd", x"4060ac2c", x"55077f3e", x"d1060001", x"55116b00", x"37a80000", x"69500000", x"ded70c95", x"5ac1cc5a", x"e00b7a41", x"80dd801b"),
	(x"66430003", x"9c2ff900", x"45aa0000", x"4c490000", x"d7e96115", x"28a308a9", x"d5c3e757", x"e14c7fae", x"2f240001", x"f2496e00", x"12790000", x"9e300000", x"57e6744f", x"4515343a", x"aedbd954", x"21fe7f84"),
	(x"69360003", x"c156e200", x"ecf20000", x"293a0000", x"513f5c55", x"afaeb14e", x"7e28bf9f", x"eed69f40", x"664e0001", x"1e197600", x"a96a0000", x"f9920000", x"7a805079", x"738484f8", x"2dc4349f", x"4a868bcb"),
	(x"65440003", x"88b3ed00", x"ae8b0000", x"75d00000", x"62956c4f", x"ba2c945a", x"eb8bf4e4", x"5a9d9fd0", x"986c0001", x"b9417300", x"8cbb0000", x"0ef20000", x"f3b128a3", x"6c507c98", x"6314978a", x"eba57454"),
	(x"97140003", x"660ee700", x"c9230000", x"de5a0000", x"d80e248f", x"b07a492e", x"30f81c8a", x"4ff560df", x"941e0001", x"f0a47c00", x"cec20000", x"52180000", x"c01b18b9", x"79d2598c", x"f6b7dcf1", x"5fee74c4"),
	(x"9b660003", x"2febe800", x"8b5a0000", x"82b00000", x"eba41495", x"a5f86c3a", x"a55b57f1", x"fbbe604f", x"6a3c0001", x"57fc7900", x"eb130000", x"a5780000", x"492a6063", x"6606a1ec", x"b8677fe4", x"fecd8b5b"),
	(x"2c2e0003", x"64e3f500", x"15980000", x"12720000", x"4ff34879", x"8cbd2498", x"6894192f", x"31e56b9f", x"de730001", x"08687000", x"9ef00000", x"0c230000", x"580131d5", x"ddcc75bd", x"4be02289", x"8f4760f5"),
	(x"205c0003", x"2d06fa00", x"57e10000", x"4e980000", x"7c597863", x"993f018c", x"fd375254", x"85ae6b0f", x"20510001", x"af307500", x"bb210000", x"fb430000", x"d130490f", x"c2188ddd", x"0530819c", x"2e649f6a"),
	(x"d20c0003", x"c3bbf000", x"30490000", x"e5120000", x"c6c230a3", x"9369dcf8", x"2644ba3a", x"90c69400", x"2c230001", x"e6d57a00", x"f9580000", x"a7a90000", x"e29a7915", x"d79aa8c9", x"9093cae7", x"9a2f9ffa"),
	(x"de7e0003", x"8a5eff00", x"72300000", x"b9f80000", x"f56800b9", x"86ebf9ec", x"b3e7f141", x"248d9490", x"d2010001", x"418d7f00", x"dc890000", x"50c90000", x"6bab01cf", x"c84e50a9", x"de4369f2", x"3b0c6065"),
	(x"eecf0001", x"6f564000", x"f33e0000", x"a79e0000", x"bdb57219", x"b711ebc5", x"4a3b40ba", x"feabf254", x"9b060002", x"61468000", x"221e0000", x"1d740000", x"36715d27", x"30495c92", x"f11336a7", x"fe1cdc7f"),
	(x"e2bd0001", x"26b34f00", x"b1470000", x"fb740000", x"8e1f4203", x"a293ced1", x"df980bc1", x"4ae0f2c4", x"65240002", x"c61e8500", x"07cf0000", x"ea140000", x"bf4025fd", x"2f9da4f2", x"bfc395b2", x"5f3f23e0"),
	(x"10ed0001", x"c80e4500", x"d6ef0000", x"50fe0000", x"34840ac3", x"a8c513a5", x"04ebe3af", x"5f880dcb", x"69560002", x"8ffb8a00", x"45b60000", x"b6fe0000", x"8cea15e7", x"3a1f81e6", x"2a60dec9", x"eb742370"),
	(x"1c9f0001", x"81eb4a00", x"94960000", x"0c140000", x"072e3ad9", x"bd4736b1", x"9148a8d4", x"ebc30d5b", x"97740002", x"28a38f00", x"60670000", x"419e0000", x"05db6d3d", x"25cb7986", x"64b07ddc", x"4a57dcef"),
	(x"abd70001", x"cae35700", x"0a540000", x"9cd60000", x"a3796635", x"94027e13", x"5c87e60a", x"2198068b", x"233b0002", x"77378600", x"15840000", x"e8c50000", x"14f03c8b", x"9e01add7", x"973720b1", x"3bdd3741"),
	(x"a7a50001", x"83065800", x"482d0000", x"c03c0000", x"90d3562f", x"81805b07", x"c924ad71", x"95d3061b", x"dd190002", x"d06f8300", x"30550000", x"1fa50000", x"9dc14451", x"81d555b7", x"d9e783a4", x"9afec8de"),
	(x"55f50001", x"6dbb5200", x"2f850000", x"6bb60000", x"2a481eef", x"8bd68673", x"1257451f", x"80bbf914", x"d16b0002", x"998a8c00", x"722c0000", x"434f0000", x"ae6b744b", x"945770a3", x"4c44c8df", x"2eb5c84e"),
	(x"59870001", x"245e5d00", x"6dfc0000", x"375c0000", x"19e22ef5", x"9e54a367", x"87f40e64", x"34f0f984", x"2f490002", x"3ed28900", x"57fd0000", x"b42f0000", x"275a0c91", x"8b8388c3", x"02946bca", x"8f9637d1"),
	(x"56f20001", x"79274600", x"c4a40000", x"522f0000", x"9f3413b5", x"19591a80", x"2c1f56ac", x"3b6a196a", x"66230002", x"d2829100", x"ecee0000", x"d38d0000", x"0a3c28a7", x"bd123801", x"818b8601", x"e4eec39e"),
	(x"5a800001", x"30c24900", x"86dd0000", x"0ec50000", x"ac9e23af", x"0cdb3f94", x"b9bc1dd7", x"8f2119fa", x"98010002", x"75da9400", x"c93f0000", x"24ed0000", x"830d507d", x"a2c6c061", x"cf5b2514", x"45cd3c01"),
	(x"a8d00001", x"de7f4300", x"e1750000", x"a54f0000", x"16056b6f", x"068de2e0", x"62cff5b9", x"9a49e6f5", x"94730002", x"3c3f9b00", x"8b460000", x"78070000", x"b0a76067", x"b744e575", x"5af86e6f", x"f1863c91"),
	(x"a4a20001", x"979a4c00", x"a30c0000", x"f9a50000", x"25af5b75", x"130fc7f4", x"f76cbec2", x"2e02e665", x"6a510002", x"9b679e00", x"ae970000", x"8f670000", x"399618bd", x"a8901d15", x"1428cd7a", x"50a5c30e"),
	(x"13ea0001", x"dc925100", x"3dce0000", x"69670000", x"81f80799", x"3a4a8f56", x"3aa3f01c", x"e459edb5", x"de1e0002", x"c4f39700", x"db740000", x"263c0000", x"28bd490b", x"135ac944", x"e7af9017", x"212f28a0"),
	(x"1f980001", x"95775e00", x"7fb70000", x"358d0000", x"b2523783", x"2fc8aa42", x"af00bb67", x"5012ed25", x"203c0002", x"63ab9200", x"fea50000", x"d15c0000", x"a18c31d1", x"0c8e3124", x"a97f3302", x"800cd73f"),
	(x"edc80001", x"7bca5400", x"181f0000", x"9e070000", x"08c97f43", x"259e7736", x"74735309", x"457a122a", x"2c4e0002", x"2a4e9d00", x"bcdc0000", x"8db60000", x"922601cb", x"190c1430", x"3cdc7879", x"3447d7af"),
	(x"e1ba0001", x"322f5b00", x"5a660000", x"c2ed0000", x"3b634f59", x"301c5222", x"e1d01872", x"f13112ba", x"d26c0002", x"8d169800", x"990d0000", x"7ad60000", x"1b177911", x"06d8ec50", x"720cdb6c", x"95642830"),
	(x"9b6b0001", x"addd6700", x"679a0000", x"376b0000", x"46cd25f9", x"fedfe06b", x"5d5c8439", x"5074942a", x"4a600002", x"7afa8300", x"bcf20000", x"ebe00000", x"35731800", x"ff39a060", x"45502db0", x"7b63e054"),
	(x"97190001", x"e4386800", x"25e30000", x"6b810000", x"756715e3", x"eb5dc57f", x"c8ffcf42", x"e43f94ba", x"b4420002", x"dda28600", x"99230000", x"1c800000", x"bc4260da", x"e0ed5800", x"0b808ea5", x"da401fcb"),
	(x"65490001", x"0a856200", x"424b0000", x"c00b0000", x"cffc5d23", x"e10b180b", x"138c272c", x"f1576bb5", x"b8300002", x"94478900", x"db5a0000", x"406a0000", x"8fe850c0", x"f56f7d14", x"9e23c5de", x"6e0b1f5b"),
	(x"693b0001", x"43606d00", x"00320000", x"9ce10000", x"fc566d39", x"f4893d1f", x"862f6c57", x"451c6b25", x"46120002", x"331f8c00", x"fe8b0000", x"b70a0000", x"06d9281a", x"eabb8574", x"d0f366cb", x"cf28e0c4"),
	(x"de730001", x"08687000", x"9ef00000", x"0c230000", x"580131d5", x"ddcc75bd", x"4be02289", x"8f4760f5", x"f25d0002", x"6c8b8500", x"8b680000", x"1e510000", x"17f279ac", x"51715125", x"23743ba6", x"bea20b6a"),
	(x"d2010001", x"418d7f00", x"dc890000", x"50c90000", x"6bab01cf", x"c84e50a9", x"de4369f2", x"3b0c6065", x"0c7f0002", x"cbd38000", x"aeb90000", x"e9310000", x"9ec30176", x"4ea5a945", x"6da498b3", x"1f81f4f5"),
	(x"20510001", x"af307500", x"bb210000", x"fb430000", x"d130490f", x"c2188ddd", x"0530819c", x"2e649f6a", x"000d0002", x"82368f00", x"ecc00000", x"b5db0000", x"ad69316c", x"5b278c51", x"f807d3c8", x"abcaf465"),
	(x"2c230001", x"e6d57a00", x"f9580000", x"a7a90000", x"e29a7915", x"d79aa8c9", x"9093cae7", x"9a2f9ffa", x"fe2f0002", x"256e8a00", x"c9110000", x"42bb0000", x"245849b6", x"44f37431", x"b6d770dd", x"0ae90bfa"),
	(x"23560001", x"bbac6100", x"50000000", x"c2da0000", x"644c4455", x"5097112e", x"3b78922f", x"95b57f14", x"b7450002", x"c93e9200", x"72020000", x"25190000", x"093e6d80", x"7262c4f3", x"35c89d16", x"6191ffb5"),
	(x"2f240001", x"f2496e00", x"12790000", x"9e300000", x"57e6744f", x"4515343a", x"aedbd954", x"21fe7f84", x"49670002", x"6e669700", x"57d30000", x"d2790000", x"800f155a", x"6db63c93", x"7b183e03", x"c0b2002a"),
	(x"dd740001", x"1cf46400", x"75d10000", x"35ba0000", x"ed7d3c8f", x"4f43e94e", x"75a8313a", x"3496808b", x"45150002", x"27839800", x"15aa0000", x"8e930000", x"b3a52540", x"78341987", x"eebb7578", x"74f900ba"),
	(x"d1060001", x"55116b00", x"37a80000", x"69500000", x"ded70c95", x"5ac1cc5a", x"e00b7a41", x"80dd801b", x"bb370002", x"80db9d00", x"307b0000", x"79f30000", x"3a945d9a", x"67e0e1e7", x"a06bd66d", x"d5daff25"),
	(x"664e0001", x"1e197600", x"a96a0000", x"f9920000", x"7a805079", x"738484f8", x"2dc4349f", x"4a868bcb", x"0f780002", x"df4f9400", x"45980000", x"d0a80000", x"2bbf0c2c", x"dc2a35b6", x"53ec8b00", x"a450148b"),
	(x"6a3c0001", x"57fc7900", x"eb130000", x"a5780000", x"492a6063", x"6606a1ec", x"b8677fe4", x"fecd8b5b", x"f15a0002", x"78179100", x"60490000", x"27c80000", x"a28e74f6", x"c3fecdd6", x"1d3c2815", x"0573eb14"),
	(x"986c0001", x"b9417300", x"8cbb0000", x"0ef20000", x"f3b128a3", x"6c507c98", x"6314978a", x"eba57454", x"fd280002", x"31f29e00", x"22300000", x"7b220000", x"912444ec", x"d67ce8c2", x"889f636e", x"b138eb84"),
	(x"941e0001", x"f0a47c00", x"cec20000", x"52180000", x"c01b18b9", x"79d2598c", x"f6b7dcf1", x"5fee74c4", x"030a0002", x"96aa9b00", x"07e10000", x"8c420000", x"18153c36", x"c9a810a2", x"c64fc07b", x"101b141b"),
	(x"3fa90001", x"74ea4300", x"6dd20000", x"510a0000", x"beb7373e", x"78611737", x"fe785bad", x"7bd4ce7f", x"3fc40002", x"b871a400", x"28560000", x"7b150000", x"ce0b4fe0", x"b6f7abce", x"5237e933", x"d5bc862a"),
	(x"33db0001", x"3d0f4c00", x"2fab0000", x"0de00000", x"8d1d0724", x"6de33223", x"6bdb10d6", x"cf9fceef", x"c1e60002", x"1f29a100", x"0d870000", x"8c750000", x"473a373a", x"a92353ae", x"1ce74a26", x"749f79b5"),
	(x"c18b0001", x"d3b24600", x"48030000", x"a66a0000", x"37864fe4", x"67b5ef57", x"b0a8f8b8", x"daf731e0", x"cd940002", x"56ccae00", x"4ffe0000", x"d09f0000", x"74900720", x"bca176ba", x"8944015d", x"c0d47925"),
	(x"cdf90001", x"9a574900", x"0a7a0000", x"fa800000", x"042c7ffe", x"7237ca43", x"250bb3c3", x"6ebc3170", x"33b60002", x"f194ab00", x"6a2f0000", x"27ff0000", x"fda17ffa", x"a3758eda", x"c794a248", x"61f786ba"),
	(x"7ab10001", x"d15f5400", x"94b80000", x"6a420000", x"a07b2312", x"5b7282e1", x"e8c4fd1d", x"a4e73aa0", x"87f90002", x"ae00a200", x"1fcc0000", x"8ea40000", x"ec8a2e4c", x"18bf5a8b", x"3413ff25", x"107d6d14"),
	(x"76c30001", x"98ba5b00", x"d6c10000", x"36a80000", x"93d11308", x"4ef0a7f5", x"7d67b666", x"10ac3a30", x"79db0002", x"0958a700", x"3a1d0000", x"79c40000", x"65bb5696", x"076ba2eb", x"7ac35c30", x"b15e928b"),
	(x"84930001", x"76075100", x"b1690000", x"9d220000", x"294a5bc8", x"44a67a81", x"a6145e08", x"05c4c53f", x"75a90002", x"40bda800", x"78640000", x"252e0000", x"5611668c", x"12e987ff", x"ef60174b", x"0515921b"),
	(x"88e10001", x"3fe25e00", x"f3100000", x"c1c80000", x"1ae06bd2", x"51245f95", x"33b71573", x"b18fc5af", x"8b8b0002", x"e7e5ad00", x"5db50000", x"d24e0000", x"df201e56", x"0d3d7f9f", x"a1b0b45e", x"a4366d84"),
	(x"87940001", x"629b4500", x"5a480000", x"a4bb0000", x"9c365692", x"d629e672", x"985c4dbb", x"be152541", x"c2e10002", x"0bb5b500", x"e6a60000", x"b5ec0000", x"f2463a60", x"3baccf5d", x"22af5995", x"cf4e99cb"),
	(x"8be60001", x"2b7e4a00", x"18310000", x"f8510000", x"af9c6688", x"c3abc366", x"0dff06c0", x"0a5e25d1", x"3cc30002", x"acedb000", x"c3770000", x"428c0000", x"7b7742ba", x"2478373d", x"6c7ffa80", x"6e6d6654"),
	(x"79b60001", x"c5c34000", x"7f990000", x"53db0000", x"15072e48", x"c9fd1e12", x"d68ceeae", x"1f36dade", x"30b10002", x"e508bf00", x"810e0000", x"1e660000", x"48dd72a0", x"31fa1229", x"f9dcb1fb", x"da2666c4"),
	(x"75c40001", x"8c264f00", x"3de00000", x"0f310000", x"26ad1e52", x"dc7f3b06", x"432fa5d5", x"ab7dda4e", x"ce930002", x"4250ba00", x"a4df0000", x"e9060000", x"c1ec0a7a", x"2e2eea49", x"b70c12ee", x"7b05995b"),
	(x"c28c0001", x"c72e5200", x"a3220000", x"9ff30000", x"82fa42be", x"f53a73a4", x"8ee0eb0b", x"6126d19e", x"7adc0002", x"1dc4b300", x"d13c0000", x"405d0000", x"d0c75bcc", x"95e43e18", x"448b4f83", x"0a8f72f5"),
	(x"cefe0001", x"8ecb5d00", x"e15b0000", x"c3190000", x"b15072a4", x"e0b856b0", x"1b43a070", x"d56dd10e", x"84fe0002", x"ba9cb600", x"f4ed0000", x"b73d0000", x"59f62316", x"8a30c678", x"0a5bec96", x"abac8d6a"),
	(x"3cae0001", x"60765700", x"86f30000", x"68930000", x"0bcb3a64", x"eaee8bc4", x"c030481e", x"c0052e01", x"888c0002", x"f379b900", x"b6940000", x"ebd70000", x"6a5c130c", x"9fb2e36c", x"9ff8a7ed", x"1fe78dfa"),
	(x"30dc0001", x"29935800", x"c48a0000", x"34790000", x"38610a7e", x"ff6caed0", x"55930365", x"744e2e91", x"76ae0002", x"5421bc00", x"93450000", x"1cb70000", x"e36d6bd6", x"80661b0c", x"d12804f8", x"bec47265"),
	(x"4a0d0001", x"b6616400", x"f9760000", x"c1ff0000", x"45cf60de", x"31af1c99", x"e91f9f2e", x"d50ba801", x"eea20002", x"a3cda700", x"b6ba0000", x"8d810000", x"cd090ac7", x"7987573c", x"e674f224", x"50c3ba01"),
	(x"467f0001", x"ff846b00", x"bb0f0000", x"9d150000", x"766550c4", x"242d398d", x"7cbcd455", x"6140a891", x"10800002", x"0495a200", x"936b0000", x"7ae10000", x"4438721d", x"6653af5c", x"a8a45131", x"f1e0459e"),
	(x"b42f0001", x"11396100", x"dca70000", x"369f0000", x"ccfe1804", x"2e7be4f9", x"a7cf3c3b", x"7428579e", x"1cf20002", x"4d70ad00", x"d1120000", x"260b0000", x"77924207", x"73d18a48", x"3d071a4a", x"45ab450e"),
	(x"b85d0001", x"58dc6e00", x"9ede0000", x"6a750000", x"ff54281e", x"3bf9c1ed", x"326c7740", x"c063570e", x"e2d00002", x"ea28a800", x"f4c30000", x"d16b0000", x"fea33add", x"6c057228", x"73d7b95f", x"e488ba91"),
	(x"0f150001", x"13d47300", x"001c0000", x"fab70000", x"5b0374f2", x"12bc894f", x"ffa3399e", x"0a385cde", x"569f0002", x"b5bca100", x"81200000", x"78300000", x"ef886b6b", x"d7cfa679", x"8050e432", x"9502513f"),
	(x"03670001", x"5a317c00", x"42650000", x"a65d0000", x"68a944e8", x"073eac5b", x"6a0072e5", x"be735c4e", x"a8bd0002", x"12e4a400", x"a4f10000", x"8f500000", x"66b913b1", x"c81b5e19", x"ce804727", x"3421aea0"),
	(x"f1370001", x"b48c7600", x"25cd0000", x"0dd70000", x"d2320c28", x"0d68712f", x"b1739a8b", x"ab1ba341", x"a4cf0002", x"5b01ab00", x"e6880000", x"d3ba0000", x"551323ab", x"dd997b0d", x"5b230c5c", x"806aae30"),
	(x"fd450001", x"fd697900", x"67b40000", x"513d0000", x"e1983c32", x"18ea543b", x"24d0d1f0", x"1f50a3d1", x"5aed0002", x"fc59ae00", x"c3590000", x"24da0000", x"dc225b71", x"c24d836d", x"15f3af49", x"214951af"),
	(x"f2300001", x"a0106200", x"ceec0000", x"344e0000", x"674e0172", x"9fe7eddc", x"8f3b8938", x"10ca433f", x"13870002", x"1009b600", x"784a0000", x"43780000", x"f1447f47", x"f4dc33af", x"96ec4282", x"4a31a5e0"),
	(x"fe420001", x"e9f56d00", x"8c950000", x"68a40000", x"54e43168", x"8a65c8c8", x"1a98c243", x"a48143af", x"eda50002", x"b751b300", x"5d9b0000", x"b4180000", x"7875079d", x"eb08cbcf", x"d83ce197", x"eb125a7f"),
	(x"0c120001", x"07486700", x"eb3d0000", x"c32e0000", x"ee7f79a8", x"803315bc", x"c1eb2a2d", x"b1e9bca0", x"e1d70002", x"feb4bc00", x"1fe20000", x"e8f20000", x"4bdf3787", x"fe8aeedb", x"4d9faaec", x"5f595aef"),
	(x"00600001", x"4ead6800", x"a9440000", x"9fc40000", x"ddd549b2", x"95b130a8", x"54486156", x"05a2bc30", x"1ff50002", x"59ecb900", x"3a330000", x"1f920000", x"c2ee4f5d", x"e15e16bb", x"034f09f9", x"fe7aa570"),
	(x"b7280001", x"05a57500", x"37860000", x"0f060000", x"7982155e", x"bcf4780a", x"99872f88", x"cff9b7e0", x"abba0002", x"0678b000", x"4fd00000", x"b6c90000", x"d3c51eeb", x"5a94c2ea", x"f0c85494", x"8ff04ede"),
	(x"bb5a0001", x"4c407a00", x"75ff0000", x"53ec0000", x"4a282544", x"a9765d1e", x"0c2464f3", x"7bb2b770", x"55980002", x"a120b500", x"6a010000", x"41a90000", x"5af46631", x"45403a8a", x"be18f781", x"2ed3b141"),
	(x"490a0001", x"a2fd7000", x"12570000", x"f8660000", x"f0b36d84", x"a320806a", x"d7578c9d", x"6eda487f", x"59ea0002", x"e8c5ba00", x"28780000", x"1d430000", x"695e562b", x"50c21f9e", x"2bbbbcfa", x"9a98b1d1"),
	(x"45780001", x"eb187f00", x"502e0000", x"a48c0000", x"c3195d9e", x"b6a2a57e", x"42f4c7e6", x"da9148ef", x"a7c80002", x"4f9dbf00", x"0da90000", x"ea230000", x"e06f2ef1", x"4f16e7fe", x"656b1fef", x"3bbb4e4e"),
	(x"9b060002", x"61468000", x"221e0000", x"1d740000", x"36715d27", x"30495c92", x"f11336a7", x"fe1cdc7f", x"75c90003", x"0e10c000", x"d1200000", x"baea0000", x"8bc42f3e", x"8758b757", x"bb28761d", x"00b72e2b"),
	(x"97740002", x"28a38f00", x"60670000", x"419e0000", x"05db6d3d", x"25cb7986", x"64b07ddc", x"4a57dcef", x"8beb0003", x"a948c500", x"f4f10000", x"4d8a0000", x"02f557e4", x"988c4f37", x"f5f8d508", x"a194d1b4"),
	(x"65240002", x"c61e8500", x"07cf0000", x"ea140000", x"bf4025fd", x"2f9da4f2", x"bfc395b2", x"5f3f23e0", x"87990003", x"e0adca00", x"b6880000", x"11600000", x"315f67fe", x"8d0e6a23", x"605b9e73", x"15dfd124"),
	(x"69560002", x"8ffb8a00", x"45b60000", x"b6fe0000", x"8cea15e7", x"3a1f81e6", x"2a60dec9", x"eb742370", x"79bb0003", x"47f5cf00", x"93590000", x"e6000000", x"b86e1f24", x"92da9243", x"2e8b3d66", x"b4fc2ebb"),
	(x"de1e0002", x"c4f39700", x"db740000", x"263c0000", x"28bd490b", x"135ac944", x"e7af9017", x"212f28a0", x"cdf40003", x"1861c600", x"e6ba0000", x"4f5b0000", x"a9454e92", x"29104612", x"dd0c600b", x"c576c515"),
	(x"d26c0002", x"8d169800", x"990d0000", x"7ad60000", x"1b177911", x"06d8ec50", x"720cdb6c", x"95642830", x"33d60003", x"bf39c300", x"c36b0000", x"b83b0000", x"20743648", x"36c4be72", x"93dcc31e", x"64553a8a"),
	(x"203c0002", x"63ab9200", x"fea50000", x"d15c0000", x"a18c31d1", x"0c8e3124", x"a97f3302", x"800cd73f", x"3fa40003", x"f6dccc00", x"81120000", x"e4d10000", x"13de0652", x"23469b66", x"067f8865", x"d01e3a1a"),
	(x"2c4e0002", x"2a4e9d00", x"bcdc0000", x"8db60000", x"922601cb", x"190c1430", x"3cdc7879", x"3447d7af", x"c1860003", x"5184c900", x"a4c30000", x"13b10000", x"9aef7e88", x"3c926306", x"48af2b70", x"713dc585"),
	(x"233b0002", x"77378600", x"15840000", x"e8c50000", x"14f03c8b", x"9e01add7", x"973720b1", x"3bdd3741", x"88ec0003", x"bdd4d100", x"1fd00000", x"74130000", x"b7895abe", x"0a03d3c4", x"cbb0c6bb", x"1a4531ca"),
	(x"2f490002", x"3ed28900", x"57fd0000", x"b42f0000", x"275a0c91", x"8b8388c3", x"02946bca", x"8f9637d1", x"76ce0003", x"1a8cd400", x"3a010000", x"83730000", x"3eb82264", x"15d72ba4", x"856065ae", x"bb66ce55"),
	(x"dd190002", x"d06f8300", x"30550000", x"1fa50000", x"9dc14451", x"81d555b7", x"d9e783a4", x"9afec8de", x"7abc0003", x"5369db00", x"78780000", x"df990000", x"0d12127e", x"00550eb0", x"10c32ed5", x"0f2dcec5"),
	(x"d16b0002", x"998a8c00", x"722c0000", x"434f0000", x"ae6b744b", x"945770a3", x"4c44c8df", x"2eb5c84e", x"849e0003", x"f431de00", x"5da90000", x"28f90000", x"84236aa4", x"1f81f6d0", x"5e138dc0", x"ae0e315a"),
	(x"66230002", x"d2829100", x"ecee0000", x"d38d0000", x"0a3c28a7", x"bd123801", x"818b8601", x"e4eec39e", x"30d10003", x"aba5d700", x"284a0000", x"81a20000", x"95083b12", x"a44b2281", x"ad94d0ad", x"df84daf4"),
	(x"6a510002", x"9b679e00", x"ae970000", x"8f670000", x"399618bd", x"a8901d15", x"1428cd7a", x"50a5c30e", x"cef30003", x"0cfdd200", x"0d9b0000", x"76c20000", x"1c3943c8", x"bb9fdae1", x"e34473b8", x"7ea7256b"),
	(x"98010002", x"75da9400", x"c93f0000", x"24ed0000", x"830d507d", x"a2c6c061", x"cf5b2514", x"45cd3c01", x"c2810003", x"4518dd00", x"4fe20000", x"2a280000", x"2f9373d2", x"ae1dfff5", x"76e738c3", x"caec25fb"),
	(x"94730002", x"3c3f9b00", x"8b460000", x"78070000", x"b0a76067", x"b744e575", x"5af86e6f", x"f1863c91", x"3ca30003", x"e240d800", x"6a330000", x"dd480000", x"a6a20b08", x"b1c90795", x"38379bd6", x"6bcfda64"),
	(x"eea20002", x"a3cda700", x"b6ba0000", x"8d810000", x"cd090ac7", x"7987573c", x"e674f224", x"50c3ba01", x"a4af0003", x"15acc300", x"4fcc0000", x"4c7e0000", x"88c66a19", x"48284ba5", x"0f6b6d0a", x"85c81200"),
	(x"e2d00002", x"ea28a800", x"f4c30000", x"d16b0000", x"fea33add", x"6c057228", x"73d7b95f", x"e488ba91", x"5a8d0003", x"b2f4c600", x"6a1d0000", x"bb1e0000", x"01f712c3", x"57fcb3c5", x"41bbce1f", x"24ebed9f"),
	(x"10800002", x"0495a200", x"936b0000", x"7ae10000", x"4438721d", x"6653af5c", x"a8a45131", x"f1e0459e", x"56ff0003", x"fb11c900", x"28640000", x"e7f40000", x"325d22d9", x"427e96d1", x"d4188564", x"90a0ed0f"),
	(x"1cf20002", x"4d70ad00", x"d1120000", x"260b0000", x"77924207", x"73d18a48", x"3d071a4a", x"45ab450e", x"a8dd0003", x"5c49cc00", x"0db50000", x"10940000", x"bb6c5a03", x"5daa6eb1", x"9ac82671", x"31831290"),
	(x"abba0002", x"0678b000", x"4fd00000", x"b6c90000", x"d3c51eeb", x"5a94c2ea", x"f0c85494", x"8ff04ede", x"1c920003", x"03ddc500", x"78560000", x"b9cf0000", x"aa470bb5", x"e660bae0", x"694f7b1c", x"4009f93e"),
	(x"a7c80002", x"4f9dbf00", x"0da90000", x"ea230000", x"e06f2ef1", x"4f16e7fe", x"656b1fef", x"3bbb4e4e", x"e2b00003", x"a485c000", x"5d870000", x"4eaf0000", x"2376736f", x"f9b44280", x"279fd809", x"e12a06a1"),
	(x"55980002", x"a120b500", x"6a010000", x"41a90000", x"5af46631", x"45403a8a", x"be18f781", x"2ed3b141", x"eec20003", x"ed60cf00", x"1ffe0000", x"12450000", x"10dc4375", x"ec366794", x"b23c9372", x"55610631"),
	(x"59ea0002", x"e8c5ba00", x"28780000", x"1d430000", x"695e562b", x"50c21f9e", x"2bbbbcfa", x"9a98b1d1", x"10e00003", x"4a38ca00", x"3a2f0000", x"e5250000", x"99ed3baf", x"f3e29ff4", x"fcec3067", x"f442f9ae"),
	(x"569f0002", x"b5bca100", x"81200000", x"78300000", x"ef886b6b", x"d7cfa679", x"8050e432", x"9502513f", x"598a0003", x"a668d200", x"813c0000", x"82870000", x"b48b1f99", x"c5732f36", x"7ff3ddac", x"9f3a0de1"),
	(x"5aed0002", x"fc59ae00", x"c3590000", x"24da0000", x"dc225b71", x"c24d836d", x"15f3af49", x"214951af", x"a7a80003", x"0130d700", x"a4ed0000", x"75e70000", x"3dba6743", x"daa7d756", x"31237eb9", x"3e19f27e"),
	(x"a8bd0002", x"12e4a400", x"a4f10000", x"8f500000", x"66b913b1", x"c81b5e19", x"ce804727", x"3421aea0", x"abda0003", x"48d5d800", x"e6940000", x"290d0000", x"0e105759", x"cf25f242", x"a48035c2", x"8a52f2ee"),
	(x"a4cf0002", x"5b01ab00", x"e6880000", x"d3ba0000", x"551323ab", x"dd997b0d", x"5b230c5c", x"806aae30", x"55f80003", x"ef8ddd00", x"c3450000", x"de6d0000", x"87212f83", x"d0f10a22", x"ea5096d7", x"2b710d71"),
	(x"13870002", x"1009b600", x"784a0000", x"43780000", x"f1447f47", x"f4dc33af", x"96ec4282", x"4a31a5e0", x"e1b70003", x"b019d400", x"b6a60000", x"77360000", x"960a7e35", x"6b3bde73", x"19d7cbba", x"5afbe6df"),
	(x"1ff50002", x"59ecb900", x"3a330000", x"1f920000", x"c2ee4f5d", x"e15e16bb", x"034f09f9", x"fe7aa570", x"1f950003", x"1741d100", x"93770000", x"80560000", x"1f3b06ef", x"74ef2613", x"570768af", x"fbd81940"),
	(x"eda50002", x"b751b300", x"5d9b0000", x"b4180000", x"7875079d", x"eb08cbcf", x"d83ce197", x"eb125a7f", x"13e70003", x"5ea4de00", x"d10e0000", x"dcbc0000", x"2c9136f5", x"616d0307", x"c2a423d4", x"4f9319d0"),
	(x"e1d70002", x"feb4bc00", x"1fe20000", x"e8f20000", x"4bdf3787", x"fe8aeedb", x"4d9faaec", x"5f595aef", x"edc50003", x"f9fcdb00", x"f4df0000", x"2bdc0000", x"a5a04e2f", x"7eb9fb67", x"8c7480c1", x"eeb0e64f"),
	(x"4a600002", x"7afa8300", x"bcf20000", x"ebe00000", x"35731800", x"ff39a060", x"45502db0", x"7b63e054", x"d10b0003", x"d727e400", x"db680000", x"dc8b0000", x"73be3df9", x"01e6400b", x"180ca989", x"2b17747e"),
	(x"46120002", x"331f8c00", x"fe8b0000", x"b70a0000", x"06d9281a", x"eabb8574", x"d0f366cb", x"cf28e0c4", x"2f290003", x"707fe100", x"feb90000", x"2beb0000", x"fa8f4523", x"1e32b86b", x"56dc0a9c", x"8a348be1"),
	(x"b4420002", x"dda28600", x"99230000", x"1c800000", x"bc4260da", x"e0ed5800", x"0b808ea5", x"da401fcb", x"235b0003", x"399aee00", x"bcc00000", x"77010000", x"c9257539", x"0bb09d7f", x"c37f41e7", x"3e7f8b71"),
	(x"b8300002", x"94478900", x"db5a0000", x"406a0000", x"8fe850c0", x"f56f7d14", x"9e23c5de", x"6e0b1f5b", x"dd790003", x"9ec2eb00", x"99110000", x"80610000", x"40140de3", x"1464651f", x"8dafe2f2", x"9f5c74ee"),
	(x"0f780002", x"df4f9400", x"45980000", x"d0a80000", x"2bbf0c2c", x"dc2a35b6", x"53ec8b00", x"a450148b", x"69360003", x"c156e200", x"ecf20000", x"293a0000", x"513f5c55", x"afaeb14e", x"7e28bf9f", x"eed69f40"),
	(x"030a0002", x"96aa9b00", x"07e10000", x"8c420000", x"18153c36", x"c9a810a2", x"c64fc07b", x"101b141b", x"97140003", x"660ee700", x"c9230000", x"de5a0000", x"d80e248f", x"b07a492e", x"30f81c8a", x"4ff560df"),
	(x"f15a0002", x"78179100", x"60490000", x"27c80000", x"a28e74f6", x"c3fecdd6", x"1d3c2815", x"0573eb14", x"9b660003", x"2febe800", x"8b5a0000", x"82b00000", x"eba41495", x"a5f86c3a", x"a55b57f1", x"fbbe604f"),
	(x"fd280002", x"31f29e00", x"22300000", x"7b220000", x"912444ec", x"d67ce8c2", x"889f636e", x"b138eb84", x"65440003", x"88b3ed00", x"ae8b0000", x"75d00000", x"62956c4f", x"ba2c945a", x"eb8bf4e4", x"5a9d9fd0"),
	(x"f25d0002", x"6c8b8500", x"8b680000", x"1e510000", x"17f279ac", x"51715125", x"23743ba6", x"bea20b6a", x"2c2e0003", x"64e3f500", x"15980000", x"12720000", x"4ff34879", x"8cbd2498", x"6894192f", x"31e56b9f"),
	(x"fe2f0002", x"256e8a00", x"c9110000", x"42bb0000", x"245849b6", x"44f37431", x"b6d770dd", x"0ae90bfa", x"d20c0003", x"c3bbf000", x"30490000", x"e5120000", x"c6c230a3", x"9369dcf8", x"2644ba3a", x"90c69400"),
	(x"0c7f0002", x"cbd38000", x"aeb90000", x"e9310000", x"9ec30176", x"4ea5a945", x"6da498b3", x"1f81f4f5", x"de7e0003", x"8a5eff00", x"72300000", x"b9f80000", x"f56800b9", x"86ebf9ec", x"b3e7f141", x"248d9490"),
	(x"000d0002", x"82368f00", x"ecc00000", x"b5db0000", x"ad69316c", x"5b278c51", x"f807d3c8", x"abcaf465", x"205c0003", x"2d06fa00", x"57e10000", x"4e980000", x"7c597863", x"993f018c", x"fd375254", x"85ae6b0f"),
	(x"b7450002", x"c93e9200", x"72020000", x"25190000", x"093e6d80", x"7262c4f3", x"35c89d16", x"6191ffb5", x"94130003", x"7292f300", x"22020000", x"e7c30000", x"6d7229d5", x"22f5d5dd", x"0eb00f39", x"f42480a1"),
	(x"bb370002", x"80db9d00", x"307b0000", x"79f30000", x"3a945d9a", x"67e0e1e7", x"a06bd66d", x"d5daff25", x"6a310003", x"d5caf600", x"07d30000", x"10a30000", x"e443510f", x"3d212dbd", x"4060ac2c", x"55077f3e"),
	(x"49670002", x"6e669700", x"57d30000", x"d2790000", x"800f155a", x"6db63c93", x"7b183e03", x"c0b2002a", x"66430003", x"9c2ff900", x"45aa0000", x"4c490000", x"d7e96115", x"28a308a9", x"d5c3e757", x"e14c7fae"),
	(x"45150002", x"27839800", x"15aa0000", x"8e930000", x"b3a52540", x"78341987", x"eebb7578", x"74f900ba", x"98610003", x"3b77fc00", x"607b0000", x"bb290000", x"5ed819cf", x"3777f0c9", x"9b134442", x"406f8031"),
	(x"3fc40002", x"b871a400", x"28560000", x"7b150000", x"ce0b4fe0", x"b6f7abce", x"5237e933", x"d5bc862a", x"006d0003", x"cc9be700", x"45840000", x"2a1f0000", x"70bc78de", x"ce96bcf9", x"ac4fb29e", x"ae684855"),
	(x"33b60002", x"f194ab00", x"6a2f0000", x"27ff0000", x"fda17ffa", x"a3758eda", x"c794a248", x"61f786ba", x"fe4f0003", x"6bc3e200", x"60550000", x"dd7f0000", x"f98d0004", x"d1424499", x"e29f118b", x"0f4bb7ca"),
	(x"c1e60002", x"1f29a100", x"0d870000", x"8c750000", x"473a373a", x"a92353ae", x"1ce74a26", x"749f79b5", x"f23d0003", x"2226ed00", x"222c0000", x"81950000", x"ca27301e", x"c4c0618d", x"773c5af0", x"bb00b75a"),
	(x"cd940002", x"56ccae00", x"4ffe0000", x"d09f0000", x"74900720", x"bca176ba", x"8944015d", x"c0d47925", x"0c1f0003", x"857ee800", x"07fd0000", x"76f50000", x"431648c4", x"db1499ed", x"39ecf9e5", x"1a2348c5"),
	(x"7adc0002", x"1dc4b300", x"d13c0000", x"405d0000", x"d0c75bcc", x"95e43e18", x"448b4f83", x"0a8f72f5", x"b8500003", x"daeae100", x"721e0000", x"dfae0000", x"523d1972", x"60de4dbc", x"ca6ba488", x"6ba9a36b"),
	(x"76ae0002", x"5421bc00", x"93450000", x"1cb70000", x"e36d6bd6", x"80661b0c", x"d12804f8", x"bec47265", x"46720003", x"7db2e400", x"57cf0000", x"28ce0000", x"db0c61a8", x"7f0ab5dc", x"84bb079d", x"ca8a5cf4"),
	(x"84fe0002", x"ba9cb600", x"f4ed0000", x"b73d0000", x"59f62316", x"8a30c678", x"0a5bec96", x"abac8d6a", x"4a000003", x"3457eb00", x"15b60000", x"74240000", x"e8a651b2", x"6a8890c8", x"11184ce6", x"7ec15c64"),
	(x"888c0002", x"f379b900", x"b6940000", x"ebd70000", x"6a5c130c", x"9fb2e36c", x"9ff8a7ed", x"1fe78dfa", x"b4220003", x"930fee00", x"30670000", x"83440000", x"61972968", x"755c68a8", x"5fc8eff3", x"dfe2a3fb"),
	(x"87f90002", x"ae00a200", x"1fcc0000", x"8ea40000", x"ec8a2e4c", x"18bf5a8b", x"3413ff25", x"107d6d14", x"fd480003", x"7f5ff600", x"8b740000", x"e4e60000", x"4cf10d5e", x"43cdd86a", x"dcd70238", x"b49a57b4"),
	(x"8b8b0002", x"e7e5ad00", x"5db50000", x"d24e0000", x"df201e56", x"0d3d7f9f", x"a1b0b45e", x"a4366d84", x"036a0003", x"d807f300", x"aea50000", x"13860000", x"c5c07584", x"5c19200a", x"9207a12d", x"15b9a82b"),
	(x"79db0002", x"0958a700", x"3a1d0000", x"79c40000", x"65bb5696", x"076ba2eb", x"7ac35c30", x"b15e928b", x"0f180003", x"91e2fc00", x"ecdc0000", x"4f6c0000", x"f66a459e", x"499b051e", x"07a4ea56", x"a1f2a8bb"),
	(x"75a90002", x"40bda800", x"78640000", x"252e0000", x"5611668c", x"12e987ff", x"ef60174b", x"0515921b", x"f13a0003", x"36baf900", x"c90d0000", x"b80c0000", x"7f5b3d44", x"564ffd7e", x"49744943", x"00d15724"),
	(x"c2e10002", x"0bb5b500", x"e6a60000", x"b5ec0000", x"f2463a60", x"3baccf5d", x"22af5995", x"cf4e99cb", x"45750003", x"692ef000", x"bcee0000", x"11570000", x"6e706cf2", x"ed85292f", x"baf3142e", x"715bbc8a"),
	(x"ce930002", x"4250ba00", x"a4df0000", x"e9060000", x"c1ec0a7a", x"2e2eea49", x"b70c12ee", x"7b05995b", x"bb570003", x"ce76f500", x"993f0000", x"e6370000", x"e7411428", x"f251d14f", x"f423b73b", x"d0784315"),
	(x"3cc30002", x"acedb000", x"c3770000", x"428c0000", x"7b7742ba", x"2478373d", x"6c7ffa80", x"6e6d6654", x"b7250003", x"8793fa00", x"db460000", x"badd0000", x"d4eb2432", x"e7d3f45b", x"6180fc40", x"64334385"),
	(x"30b10002", x"e508bf00", x"810e0000", x"1e660000", x"48dd72a0", x"31fa1229", x"f9dcb1fb", x"da2666c4", x"49070003", x"20cbff00", x"fe970000", x"4dbd0000", x"5dda5ce8", x"f8070c3b", x"2f505f55", x"c510bc1a")
    ),(
	(x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000"),
	(x"86790000", x"3f390002", x"e19ae000", x"98560000", x"9565670e", x"4e88c8ea", x"d3dd4944", x"161ddab9", x"30b70000", x"e5d00000", x"f4f46000", x"42c40000", x"63b83d6a", x"78ba9460", x"21afa1ea", x"b0a51834"),
	(x"30b70000", x"e5d00000", x"f4f46000", x"42c40000", x"63b83d6a", x"78ba9460", x"21afa1ea", x"b0a51834", x"b6ce0000", x"dae90002", x"156e8000", x"da920000", x"f6dd5a64", x"36325c8a", x"f272e8ae", x"a6b8c28d"),
	(x"b6ce0000", x"dae90002", x"156e8000", x"da920000", x"f6dd5a64", x"36325c8a", x"f272e8ae", x"a6b8c28d", x"86790000", x"3f390002", x"e19ae000", x"98560000", x"9565670e", x"4e88c8ea", x"d3dd4944", x"161ddab9"),
	(x"14190000", x"23ca003c", x"50df0000", x"44b60000", x"1b6c67b0", x"3cf3ac75", x"61e610b0", x"dbcadb80", x"e3430000", x"3a4e0014", x"f2c60000", x"aa4e0000", x"db1e42a6", x"256bbe15", x"123db156", x"3a4e99d7"),
	(x"92600000", x"1cf3003e", x"b145e000", x"dce00000", x"8e0900be", x"727b649f", x"b23b59f4", x"cdd70139", x"d3f40000", x"df9e0014", x"06326000", x"e88a0000", x"b8a67fcc", x"5dd12a75", x"339210bc", x"8aeb81e3"),
	(x"24ae0000", x"c61a003c", x"a42b6000", x"06720000", x"78d45ada", x"44493815", x"4049b15a", x"6b6fc3b4", x"558d0000", x"e0a70016", x"e7a88000", x"70dc0000", x"2dc318c2", x"1359e29f", x"e04f59f8", x"9cf65b5a"),
	(x"a2d70000", x"f923003e", x"45b18000", x"9e240000", x"edb13dd4", x"0ac1f0ff", x"9394f81e", x"7d72190d", x"653a0000", x"05770016", x"135ce000", x"32180000", x"4e7b25a8", x"6be376ff", x"c1e0f812", x"2c53436e"),
	(x"e3430000", x"3a4e0014", x"f2c60000", x"aa4e0000", x"db1e42a6", x"256bbe15", x"123db156", x"3a4e99d7", x"f75a0000", x"19840028", x"a2190000", x"eef80000", x"c0722516", x"19981260", x"73dba1e6", x"e1844257"),
	(x"653a0000", x"05770016", x"135ce000", x"32180000", x"4e7b25a8", x"6be376ff", x"c1e0f812", x"2c53436e", x"c7ed0000", x"fc540028", x"56ed6000", x"ac3c0000", x"a3ca187c", x"61228600", x"5274000c", x"51215a63"),
	(x"d3f40000", x"df9e0014", x"06326000", x"e88a0000", x"b8a67fcc", x"5dd12a75", x"339210bc", x"8aeb81e3", x"41940000", x"c36d002a", x"b7778000", x"346a0000", x"36af7f72", x"2faa4eea", x"81a94948", x"473c80da"),
	(x"558d0000", x"e0a70016", x"e7a88000", x"70dc0000", x"2dc318c2", x"1359e29f", x"e04f59f8", x"9cf65b5a", x"71230000", x"26bd002a", x"4383e000", x"76ae0000", x"55174218", x"5710da8a", x"a006e8a2", x"f79998ee"),
	(x"f75a0000", x"19840028", x"a2190000", x"eef80000", x"c0722516", x"19981260", x"73dba1e6", x"e1844257", x"14190000", x"23ca003c", x"50df0000", x"44b60000", x"1b6c67b0", x"3cf3ac75", x"61e610b0", x"dbcadb80"),
	(x"71230000", x"26bd002a", x"4383e000", x"76ae0000", x"55174218", x"5710da8a", x"a006e8a2", x"f79998ee", x"24ae0000", x"c61a003c", x"a42b6000", x"06720000", x"78d45ada", x"44493815", x"4049b15a", x"6b6fc3b4"),
	(x"c7ed0000", x"fc540028", x"56ed6000", x"ac3c0000", x"a3ca187c", x"61228600", x"5274000c", x"51215a63", x"a2d70000", x"f923003e", x"45b18000", x"9e240000", x"edb13dd4", x"0ac1f0ff", x"9394f81e", x"7d72190d"),
	(x"41940000", x"c36d002a", x"b7778000", x"346a0000", x"36af7f72", x"2faa4eea", x"81a94948", x"473c80da", x"92600000", x"1cf3003e", x"b145e000", x"dce00000", x"8e0900be", x"727b649f", x"b23b59f4", x"cdd70139"),
	(x"54500000", x"0671005c", x"25ae0000", x"6a1e0000", x"2ea54edf", x"664e8512", x"bfba18c3", x"7e715d17", x"bc8d0000", x"fc3b0018", x"19830000", x"d10b0000", x"ae1878c4", x"42a69856", x"0012da37", x"2c3b504e"),
	(x"d2290000", x"3948005e", x"c434e000", x"f2480000", x"bbc029d1", x"28c64df8", x"6c675187", x"686c87ae", x"8c3a0000", x"19eb0018", x"ed776000", x"93cf0000", x"cda045ae", x"3a1c0c36", x"21bd7bdd", x"9c9e487a"),
	(x"64e70000", x"e3a1005c", x"d15a6000", x"28da0000", x"4d1d73b5", x"1ef41172", x"9e15b929", x"ced44523", x"0a430000", x"26d2001a", x"0ced8000", x"0b990000", x"58c522a0", x"7494c4dc", x"f2603299", x"8a8392c3"),
	(x"e29e0000", x"dc98005e", x"30c08000", x"b08c0000", x"d87814bb", x"507cd998", x"4dc8f06d", x"d8c99f9a", x"3af40000", x"c302001a", x"f819e000", x"495d0000", x"3b7d1fca", x"0c2e50bc", x"d3cf9373", x"3a268af7"),
	(x"40490000", x"25bb0060", x"75710000", x"2ea80000", x"35c9296f", x"5abd2967", x"de5c0873", x"a5bb8697", x"5fce0000", x"c675000c", x"eb450000", x"7b450000", x"75063a62", x"67cd2643", x"122f6b61", x"1675c999"),
	(x"c6300000", x"1a820062", x"94ebe000", x"b6fe0000", x"a0ac4e61", x"1435e18d", x"0d814137", x"b3a65c2e", x"6f790000", x"23a5000c", x"1fb16000", x"39810000", x"16be0708", x"1f77b223", x"3380ca8b", x"a6d0d1ad"),
	(x"70fe0000", x"c06b0060", x"81856000", x"6c6c0000", x"56711405", x"2207bd07", x"fff3a999", x"151e9ea3", x"e9000000", x"1c9c000e", x"fe2b8000", x"a1d70000", x"83db6006", x"51ff7ac9", x"e05d83cf", x"b0cd0b14"),
	(x"f6870000", x"ff520062", x"601f8000", x"f43a0000", x"c314730b", x"6c8f75ed", x"2c2ee0dd", x"0303441a", x"d9b70000", x"f94c000e", x"0adfe000", x"e3130000", x"e0635d6c", x"2945eea9", x"c1f22225", x"00681320"),
	(x"b7130000", x"3c3f0048", x"d7680000", x"c0500000", x"f5bb0c79", x"43253b07", x"ad87a995", x"443fc4c0", x"4bd70000", x"e5bf0030", x"bb9a0000", x"3ff30000", x"6e6a5dd2", x"5b3e8a36", x"73c97bd1", x"cdbf1219"),
	(x"316a0000", x"0306004a", x"36f2e000", x"58060000", x"60de6b77", x"0dadf3ed", x"7e5ae0d1", x"52221e79", x"7b600000", x"006f0030", x"4f6e6000", x"7d370000", x"0dd260b8", x"23841e56", x"5266da3b", x"7d1a0a2d"),
	(x"87a40000", x"d9ef0048", x"239c6000", x"82940000", x"96033113", x"3b9faf67", x"8c28087f", x"f49adcf4", x"fd190000", x"3f560032", x"aef48000", x"e5610000", x"98b707b6", x"6d0cd6bc", x"81bb937f", x"6b07d094"),
	(x"01dd0000", x"e6d6004a", x"c2068000", x"1ac20000", x"0366561d", x"7517678d", x"5ff5413b", x"e287064d", x"cdae0000", x"da860032", x"5a00e000", x"a7a50000", x"fb0f3adc", x"15b642dc", x"a0143295", x"dba2c8a0"),
	(x"a30a0000", x"1ff50074", x"87b70000", x"84e60000", x"eed76bc9", x"7fd69772", x"cc61b925", x"9ff51f40", x"a8940000", x"dff10024", x"495c0000", x"95bd0000", x"b5741f74", x"7e553423", x"61f4ca87", x"f7f18bce"),
	(x"25730000", x"20cc0076", x"662de000", x"1cb00000", x"7bb20cc7", x"315e5f98", x"1fbcf061", x"89e8c5f9", x"98230000", x"3a210024", x"bda86000", x"d7790000", x"d6cc221e", x"06efa043", x"405b6b6d", x"475493fa"),
	(x"93bd0000", x"fa250074", x"73436000", x"c6220000", x"8d6f56a3", x"076c0312", x"edce18cf", x"2f500774", x"1e5a0000", x"05180026", x"5c328000", x"4f2f0000", x"43a94510", x"486768a9", x"93862229", x"51494943"),
	(x"15c40000", x"c51c0076", x"92d98000", x"5e740000", x"180a31ad", x"49e4cbf8", x"3e13518b", x"394dddcd", x"2eed0000", x"e0c80026", x"a8c6e000", x"0deb0000", x"2011787a", x"30ddfcc9", x"b22983c3", x"e1ec5177"),
	(x"bc8d0000", x"fc3b0018", x"19830000", x"d10b0000", x"ae1878c4", x"42a69856", x"0012da37", x"2c3b504e", x"e8dd0000", x"fa4a0044", x"3c2d0000", x"bb150000", x"80bd361b", x"24e81d44", x"bfa8c2f4", x"524a0d59"),
	(x"3af40000", x"c302001a", x"f819e000", x"495d0000", x"3b7d1fca", x"0c2e50bc", x"d3cf9373", x"3a268af7", x"d86a0000", x"1f9a0044", x"c8d96000", x"f9d10000", x"e3050b71", x"5c528924", x"9e07631e", x"e2ef156d"),
	(x"8c3a0000", x"19eb0018", x"ed776000", x"93cf0000", x"cda045ae", x"3a1c0c36", x"21bd7bdd", x"9c9e487a", x"5e130000", x"20a30046", x"29438000", x"61870000", x"76606c7f", x"12da41ce", x"4dda2a5a", x"f4f2cfd4"),
	(x"0a430000", x"26d2001a", x"0ced8000", x"0b990000", x"58c522a0", x"7494c4dc", x"f2603299", x"8a8392c3", x"6ea40000", x"c5730046", x"ddb7e000", x"23430000", x"15d85115", x"6a60d5ae", x"6c758bb0", x"4457d7e0"),
	(x"a8940000", x"dff10024", x"495c0000", x"95bd0000", x"b5741f74", x"7e553423", x"61f4ca87", x"f7f18bce", x"0b9e0000", x"c0040050", x"ceeb0000", x"115b0000", x"5ba374bd", x"0183a351", x"ad9573a2", x"6804948e"),
	(x"2eed0000", x"e0c80026", x"a8c6e000", x"0deb0000", x"2011787a", x"30ddfcc9", x"b22983c3", x"e1ec5177", x"3b290000", x"25d40050", x"3a1f6000", x"539f0000", x"381b49d7", x"79393731", x"8c3ad248", x"d8a18cba"),
	(x"98230000", x"3a210024", x"bda86000", x"d7790000", x"d6cc221e", x"06efa043", x"405b6b6d", x"475493fa", x"bd500000", x"1aed0052", x"db858000", x"cbc90000", x"ad7e2ed9", x"37b1ffdb", x"5fe79b0c", x"cebc5603"),
	(x"1e5a0000", x"05180026", x"5c328000", x"4f2f0000", x"43a94510", x"486768a9", x"93862229", x"51494943", x"8de70000", x"ff3d0052", x"2f71e000", x"890d0000", x"cec613b3", x"4f0b6bbb", x"7e483ae6", x"7e194e37"),
	(x"5fce0000", x"c675000c", x"eb450000", x"7b450000", x"75063a62", x"67cd2643", x"122f6b61", x"1675c999", x"1f870000", x"e3ce006c", x"9e340000", x"55ed0000", x"40cf130d", x"3d700f24", x"cc736312", x"b3ce4f0e"),
	(x"d9b70000", x"f94c000e", x"0adfe000", x"e3130000", x"e0635d6c", x"2945eea9", x"c1f22225", x"00681320", x"2f300000", x"061e006c", x"6ac06000", x"17290000", x"23772e67", x"45ca9b44", x"eddcc2f8", x"036b573a"),
	(x"6f790000", x"23a5000c", x"1fb16000", x"39810000", x"16be0708", x"1f77b223", x"3380ca8b", x"a6d0d1ad", x"a9490000", x"3927006e", x"8b5a8000", x"8f7f0000", x"b6124969", x"0b4253ae", x"3e018bbc", x"15768d83"),
	(x"e9000000", x"1c9c000e", x"fe2b8000", x"a1d70000", x"83db6006", x"51ff7ac9", x"e05d83cf", x"b0cd0b14", x"99fe0000", x"dcf7006e", x"7faee000", x"cdbb0000", x"d5aa7403", x"73f8c7ce", x"1fae2a56", x"a5d395b7"),
	(x"4bd70000", x"e5bf0030", x"bb9a0000", x"3ff30000", x"6e6a5dd2", x"5b3e8a36", x"73c97bd1", x"cdbf1219", x"fcc40000", x"d9800078", x"6cf20000", x"ffa30000", x"9bd151ab", x"181bb131", x"de4ed244", x"8980d6d9"),
	(x"cdae0000", x"da860032", x"5a00e000", x"a7a50000", x"fb0f3adc", x"15b642dc", x"a0143295", x"dba2c8a0", x"cc730000", x"3c500078", x"98066000", x"bd670000", x"f8696cc1", x"60a12551", x"ffe173ae", x"3925ceed"),
	(x"7b600000", x"006f0030", x"4f6e6000", x"7d370000", x"0dd260b8", x"23841e56", x"5266da3b", x"7d1a0a2d", x"4a0a0000", x"0369007a", x"799c8000", x"25310000", x"6d0c0bcf", x"2e29edbb", x"2c3c3aea", x"2f381454"),
	(x"fd190000", x"3f560032", x"aef48000", x"e5610000", x"98b707b6", x"6d0cd6bc", x"81bb937f", x"6b07d094", x"7abd0000", x"e6b9007a", x"8d68e000", x"67f50000", x"0eb436a5", x"569379db", x"0d939b00", x"9f9d0c60"),
	(x"e8dd0000", x"fa4a0044", x"3c2d0000", x"bb150000", x"80bd361b", x"24e81d44", x"bfa8c2f4", x"524a0d59", x"54500000", x"0671005c", x"25ae0000", x"6a1e0000", x"2ea54edf", x"664e8512", x"bfba18c3", x"7e715d17"),
	(x"6ea40000", x"c5730046", x"ddb7e000", x"23430000", x"15d85115", x"6a60d5ae", x"6c758bb0", x"4457d7e0", x"64e70000", x"e3a1005c", x"d15a6000", x"28da0000", x"4d1d73b5", x"1ef41172", x"9e15b929", x"ced44523"),
	(x"d86a0000", x"1f9a0044", x"c8d96000", x"f9d10000", x"e3050b71", x"5c528924", x"9e07631e", x"e2ef156d", x"e29e0000", x"dc98005e", x"30c08000", x"b08c0000", x"d87814bb", x"507cd998", x"4dc8f06d", x"d8c99f9a"),
	(x"5e130000", x"20a30046", x"29438000", x"61870000", x"76606c7f", x"12da41ce", x"4dda2a5a", x"f4f2cfd4", x"d2290000", x"3948005e", x"c434e000", x"f2480000", x"bbc029d1", x"28c64df8", x"6c675187", x"686c87ae"),
	(x"fcc40000", x"d9800078", x"6cf20000", x"ffa30000", x"9bd151ab", x"181bb131", x"de4ed244", x"8980d6d9", x"b7130000", x"3c3f0048", x"d7680000", x"c0500000", x"f5bb0c79", x"43253b07", x"ad87a995", x"443fc4c0"),
	(x"7abd0000", x"e6b9007a", x"8d68e000", x"67f50000", x"0eb436a5", x"569379db", x"0d939b00", x"9f9d0c60", x"87a40000", x"d9ef0048", x"239c6000", x"82940000", x"96033113", x"3b9faf67", x"8c28087f", x"f49adcf4"),
	(x"cc730000", x"3c500078", x"98066000", x"bd670000", x"f8696cc1", x"60a12551", x"ffe173ae", x"3925ceed", x"01dd0000", x"e6d6004a", x"c2068000", x"1ac20000", x"0366561d", x"7517678d", x"5ff5413b", x"e287064d"),
	(x"4a0a0000", x"0369007a", x"799c8000", x"25310000", x"6d0c0bcf", x"2e29edbb", x"2c3c3aea", x"2f381454", x"316a0000", x"0306004a", x"36f2e000", x"58060000", x"60de6b77", x"0dadf3ed", x"7e5ae0d1", x"52221e79"),
	(x"0b9e0000", x"c0040050", x"ceeb0000", x"115b0000", x"5ba374bd", x"0183a351", x"ad9573a2", x"6804948e", x"a30a0000", x"1ff50074", x"87b70000", x"84e60000", x"eed76bc9", x"7fd69772", x"cc61b925", x"9ff51f40"),
	(x"8de70000", x"ff3d0052", x"2f71e000", x"890d0000", x"cec613b3", x"4f0b6bbb", x"7e483ae6", x"7e194e37", x"93bd0000", x"fa250074", x"73436000", x"c6220000", x"8d6f56a3", x"076c0312", x"edce18cf", x"2f500774"),
	(x"3b290000", x"25d40050", x"3a1f6000", x"539f0000", x"381b49d7", x"79393731", x"8c3ad248", x"d8a18cba", x"15c40000", x"c51c0076", x"92d98000", x"5e740000", x"180a31ad", x"49e4cbf8", x"3e13518b", x"394dddcd"),
	(x"bd500000", x"1aed0052", x"db858000", x"cbc90000", x"ad7e2ed9", x"37b1ffdb", x"5fe79b0c", x"cebc5603", x"25730000", x"20cc0076", x"662de000", x"1cb00000", x"7bb20cc7", x"315e5f98", x"1fbcf061", x"89e8c5f9"),
	(x"1f870000", x"e3ce006c", x"9e340000", x"55ed0000", x"40cf130d", x"3d700f24", x"cc736312", x"b3ce4f0e", x"40490000", x"25bb0060", x"75710000", x"2ea80000", x"35c9296f", x"5abd2967", x"de5c0873", x"a5bb8697"),
	(x"99fe0000", x"dcf7006e", x"7faee000", x"cdbb0000", x"d5aa7403", x"73f8c7ce", x"1fae2a56", x"a5d395b7", x"70fe0000", x"c06b0060", x"81856000", x"6c6c0000", x"56711405", x"2207bd07", x"fff3a999", x"151e9ea3"),
	(x"2f300000", x"061e006c", x"6ac06000", x"17290000", x"23772e67", x"45ca9b44", x"eddcc2f8", x"036b573a", x"f6870000", x"ff520062", x"601f8000", x"f43a0000", x"c314730b", x"6c8f75ed", x"2c2ee0dd", x"0303441a"),
	(x"a9490000", x"3927006e", x"8b5a8000", x"8f7f0000", x"b6124969", x"0b4253ae", x"3e018bbc", x"15768d83", x"c6300000", x"1a820062", x"94ebe000", x"b6fe0000", x"a0ac4e61", x"1435e18d", x"0d814137", x"b3a65c2e"),
	(x"69510000", x"d4e1009c", x"c3230000", x"ac2f0000", x"e4950bae", x"cea415dc", x"87ec287c", x"bce1a3ce", x"c6730000", x"af8d000c", x"a4c10000", x"218d0000", x"23111587", x"7913512f", x"1d28ac88", x"378dd173"),
	(x"ef280000", x"ebd8009e", x"22b9e000", x"34790000", x"71f06ca0", x"802cdd36", x"54316138", x"aafc7977", x"f6c40000", x"4a5d000c", x"50356000", x"63490000", x"40a928ed", x"01a9c54f", x"3c870d62", x"8728c947"),
	(x"59e60000", x"3131009c", x"37d76000", x"eeeb0000", x"872d36c4", x"b61e81bc", x"a6438996", x"0c44bbfa", x"70bd0000", x"7564000e", x"b1af8000", x"fb1f0000", x"d5cc4fe3", x"4f210da5", x"ef5a4426", x"913513fe"),
	(x"df9f0000", x"0e08009e", x"d64d8000", x"76bd0000", x"124851ca", x"f8964956", x"759ec0d2", x"1a596143", x"400a0000", x"90b4000e", x"455be000", x"b9db0000", x"b6747289", x"379b99c5", x"cef5e5cc", x"21900bca"),
	(x"7d480000", x"f72b00a0", x"93fc0000", x"e8990000", x"fff96c1e", x"f257b9a9", x"e60a38cc", x"672b784e", x"25300000", x"95c30018", x"56070000", x"8bc30000", x"f80f5721", x"5c78ef3a", x"0f151dde", x"0dc348a4"),
	(x"fb310000", x"c81200a2", x"7266e000", x"70cf0000", x"6a9c0b10", x"bcdf7143", x"35d77188", x"7136a2f7", x"15870000", x"70130018", x"a2f36000", x"c9070000", x"9bb76a4b", x"24c27b5a", x"2ebabc34", x"bd665090"),
	(x"4dff0000", x"12fb00a0", x"67086000", x"aa5d0000", x"9c415174", x"8aed2dc9", x"c7a59926", x"d78e607a", x"93fe0000", x"4f2a001a", x"43698000", x"51510000", x"0ed20d45", x"6a4ab3b0", x"fd67f570", x"ab7b8a29"),
	(x"cb860000", x"2dc200a2", x"86928000", x"320b0000", x"0924367a", x"c465e523", x"1478d062", x"c193bac3", x"a3490000", x"aafa001a", x"b79de000", x"13950000", x"6d6a302f", x"12f027d0", x"dcc8549a", x"1bde921d"),
	(x"8a120000", x"eeaf0088", x"31e50000", x"06610000", x"3f8b4908", x"ebcfabc9", x"95d1992a", x"86af3a19", x"31290000", x"b6090024", x"06d80000", x"cf750000", x"e3633091", x"608b434f", x"6ef30d6e", x"d6099324"),
	(x"0c6b0000", x"d196008a", x"d07fe000", x"9e370000", x"aaee2e06", x"a5476323", x"460cd06e", x"90b2e0a0", x"019e0000", x"53d90024", x"f22c6000", x"8db10000", x"80db0dfb", x"1831d72f", x"4f5cac84", x"66ac8b10"),
	(x"baa50000", x"0b7f0088", x"c5116000", x"44a50000", x"5c337462", x"93753fa9", x"b47e38c0", x"360a222d", x"87e70000", x"6ce00026", x"13b68000", x"15e70000", x"15be6af5", x"56b91fc5", x"9c81e5c0", x"70b151a9"),
	(x"3cdc0000", x"3446008a", x"248b8000", x"dcf30000", x"c956136c", x"ddfdf743", x"67a37184", x"2017f894", x"b7500000", x"89300026", x"e742e000", x"57230000", x"7606579f", x"2e038ba5", x"bd2e442a", x"c014499d"),
	(x"9e0b0000", x"cd6500b4", x"613a0000", x"42d70000", x"24e72eb8", x"d73c07bc", x"f437899a", x"5d65e199", x"d26a0000", x"8c470030", x"f41e0000", x"653b0000", x"387d7237", x"45e0fd5a", x"7ccebc38", x"ec470af3"),
	(x"18720000", x"f25c00b6", x"80a0e000", x"da810000", x"b18249b6", x"99b4cf56", x"27eac0de", x"4b783b20", x"e2dd0000", x"69970030", x"00ea6000", x"27ff0000", x"5bc54f5d", x"3d5a693a", x"5d611dd2", x"5ce212c7"),
	(x"aebc0000", x"28b500b4", x"95ce6000", x"00130000", x"475f13d2", x"af8693dc", x"d5982870", x"edc0f9ad", x"64a40000", x"56ae0032", x"e1708000", x"bfa90000", x"cea02853", x"73d2a1d0", x"8ebc5496", x"4affc87e"),
	(x"28c50000", x"178c00b6", x"74548000", x"98450000", x"d23a74dc", x"e10e5b36", x"06456134", x"fbdd2314", x"54130000", x"b37e0032", x"1584e000", x"fd6d0000", x"ad181539", x"0b6835b0", x"af13f57c", x"fa5ad04a"),
	(x"3d010000", x"d29000c0", x"e68d0000", x"c6310000", x"ca304571", x"a8ea90ce", x"385630bf", x"c290fed9", x"7afe0000", x"53b60014", x"bd420000", x"f0860000", x"8d096d43", x"3bb5c979", x"1d3a76bf", x"1bb6813d"),
	(x"bb780000", x"eda900c2", x"0717e000", x"5e670000", x"5f55227f", x"e6625824", x"eb8b79fb", x"d48d2460", x"4a490000", x"b6660014", x"49b66000", x"b2420000", x"eeb15029", x"430f5d19", x"3c95d755", x"ab139909"),
	(x"0db60000", x"374000c0", x"12796000", x"84f50000", x"a988781b", x"d05004ae", x"19f99155", x"7235e6ed", x"cc300000", x"895f0016", x"a82c8000", x"2a140000", x"7bd43727", x"0d8795f3", x"ef489e11", x"bd0e43b0"),
	(x"8bcf0000", x"087900c2", x"f3e38000", x"1ca30000", x"3ced1f15", x"9ed8cc44", x"ca24d811", x"64283c54", x"fc870000", x"6c8f0016", x"5cd8e000", x"68d00000", x"186c0a4d", x"753d0193", x"cee73ffb", x"0dab5b84"),
	(x"29180000", x"f15a00fc", x"b6520000", x"82870000", x"d15c22c1", x"94193cbb", x"59b0200f", x"195a2559", x"99bd0000", x"69f80000", x"4f840000", x"5ac80000", x"56172fe5", x"1ede776c", x"0f07c7e9", x"21f818ea"),
	(x"af610000", x"ce6300fe", x"57c8e000", x"1ad10000", x"443945cf", x"da91f451", x"8a6d694b", x"0f47ffe0", x"a90a0000", x"8c280000", x"bb706000", x"180c0000", x"35af128f", x"6664e30c", x"2ea86603", x"915d00de"),
	(x"19af0000", x"148a00fc", x"42a66000", x"c0430000", x"b2e41fab", x"eca3a8db", x"781f81e5", x"a9ff3d6d", x"2f730000", x"b3110002", x"5aea8000", x"805a0000", x"a0ca7581", x"28ec2be6", x"fd752f47", x"8740da67"),
	(x"9fd60000", x"2bb300fe", x"a33c8000", x"58150000", x"278178a5", x"a22b6031", x"abc2c8a1", x"bfe2e7d4", x"1fc40000", x"56c10002", x"ae1ee000", x"c29e0000", x"c37248eb", x"5056bf86", x"dcda8ead", x"37e5c253"),
	(x"de420000", x"e8de00d4", x"144b0000", x"6c7f0000", x"112e07d7", x"8d812edb", x"2a6b81e9", x"f8de670e", x"8da40000", x"4a32003c", x"1f5b0000", x"1e7e0000", x"4d7b4855", x"222ddb19", x"6ee1d759", x"fa32c36a"),
	(x"583b0000", x"d7e700d6", x"f5d1e000", x"f4290000", x"844b60d9", x"c309e631", x"f9b6c8ad", x"eec3bdb7", x"bd130000", x"afe2003c", x"ebaf6000", x"5cba0000", x"2ec3753f", x"5a974f79", x"4f4e76b3", x"4a97db5e"),
	(x"eef50000", x"0d0e00d4", x"e0bf6000", x"2ebb0000", x"72963abd", x"f53bbabb", x"0bc42003", x"487b7f3a", x"3b6a0000", x"90db003e", x"0a358000", x"c4ec0000", x"bba61231", x"141f8793", x"9c933ff7", x"5c8a01e7"),
	(x"688c0000", x"323700d6", x"01258000", x"b6ed0000", x"e7f35db3", x"bbb37251", x"d8196947", x"5e66a583", x"0bdd0000", x"750b003e", x"fec1e000", x"86280000", x"d81e2f5b", x"6ca513f3", x"bd3c9e1d", x"ec2f19d3"),
	(x"ca5b0000", x"cb1400e8", x"44940000", x"28c90000", x"0a426067", x"b17282ae", x"4b8d9159", x"2314bc8e", x"6ee70000", x"707c0028", x"ed9d0000", x"b4300000", x"96650af3", x"0746650c", x"7cdc660f", x"c07c5abd"),
	(x"4c220000", x"f42d00ea", x"a50ee000", x"b09f0000", x"9f270769", x"fffa4a44", x"9850d81d", x"35096637", x"5e500000", x"95ac0028", x"19696000", x"f6f40000", x"f5dd3799", x"7ffcf16c", x"5d73c7e5", x"70d94289"),
	(x"faec0000", x"2ec400e8", x"b0606000", x"6a0d0000", x"69fa5d0d", x"c9c816ce", x"6a2230b3", x"93b1a4ba", x"d8290000", x"aa95002a", x"f8f38000", x"6ea20000", x"60b85097", x"31743986", x"8eae8ea1", x"66c49830"),
	(x"7c950000", x"11fd00ea", x"51fa8000", x"f25b0000", x"fc9f3a03", x"8740de24", x"b9ff79f7", x"85ac7e03", x"e89e0000", x"4f45002a", x"0c07e000", x"2c660000", x"03006dfd", x"49ceade6", x"af012f4b", x"d6618004"),
	(x"d5dc0000", x"28da0084", x"daa00000", x"7d240000", x"4a8d736a", x"8c028d8a", x"87fef24b", x"90daf380", x"2eae0000", x"55c70048", x"98ec0000", x"9a980000", x"a3ac239c", x"5dfb4c6b", x"a2806e7c", x"65c7dc2a"),
	(x"53a50000", x"17e30086", x"3b3ae000", x"e5720000", x"dfe81464", x"c28a4560", x"5423bb0f", x"86c72939", x"1e190000", x"b0170048", x"6c186000", x"d85c0000", x"c0141ef6", x"2541d80b", x"832fcf96", x"d562c41e"),
	(x"e56b0000", x"cd0a0084", x"2e546000", x"3fe00000", x"29354e00", x"f4b819ea", x"a65153a1", x"207febb4", x"98600000", x"8f2e004a", x"8d828000", x"400a0000", x"557179f8", x"6bc910e1", x"50f286d2", x"c37f1ea7"),
	(x"63120000", x"f2330086", x"cfce8000", x"a7b60000", x"bc50290e", x"ba30d100", x"758c1ae5", x"3662310d", x"a8d70000", x"6afe004a", x"7976e000", x"02ce0000", x"36c94492", x"13738481", x"715d2738", x"73da0693"),
	(x"c1c50000", x"0b1000b8", x"8a7f0000", x"39920000", x"51e114da", x"b0f121ff", x"e618e2fb", x"4b102800", x"cded0000", x"6f89005c", x"6a2a0000", x"30d60000", x"78b2613a", x"7890f27e", x"b0bddf2a", x"5f8945fd"),
	(x"47bc0000", x"342900ba", x"6be5e000", x"a1c40000", x"c48473d4", x"fe79e915", x"35c5abbf", x"5d0df2b9", x"fd5a0000", x"8a59005c", x"9ede6000", x"72120000", x"1b0a5c50", x"002a661e", x"91127ec0", x"ef2c5dc9"),
	(x"f1720000", x"eec000b8", x"7e8b6000", x"7b560000", x"325929b0", x"c84bb59f", x"c7b74311", x"fbb53034", x"7b230000", x"b560005e", x"7f448000", x"ea440000", x"8e6f3b5e", x"4ea2aef4", x"42cf3784", x"f9318770"),
	(x"770b0000", x"d1f900ba", x"9f118000", x"e3000000", x"a73c4ebe", x"86c37d75", x"146a0a55", x"eda8ea8d", x"4b940000", x"50b0005e", x"8bb0e000", x"a8800000", x"edd70634", x"36183a94", x"6360966e", x"49949f44"),
	(x"369f0000", x"12940090", x"28660000", x"d76a0000", x"919331cc", x"a969339f", x"95c3431d", x"aa946a57", x"d9f40000", x"4c430060", x"3af50000", x"74600000", x"63de068a", x"44635e0b", x"d15bcf9a", x"84439e7d"),
	(x"b0e60000", x"2dad0092", x"c9fce000", x"4f3c0000", x"04f656c2", x"e7e1fb75", x"461e0a59", x"bc89b0ee", x"e9430000", x"a9930060", x"ce016000", x"36a40000", x"00663be0", x"3cd9ca6b", x"f0f46e70", x"34e68649"),
	(x"06280000", x"f7440090", x"dc926000", x"95ae0000", x"f22b0ca6", x"d1d3a7ff", x"b46ce2f7", x"1a317263", x"6f3a0000", x"96aa0062", x"2f9b8000", x"aef20000", x"95035cee", x"72510281", x"23292734", x"22fb5cf0"),
	(x"80510000", x"c87d0092", x"3d088000", x"0df80000", x"674e6ba8", x"9f5b6f15", x"67b1abb3", x"0c2ca8da", x"5f8d0000", x"737a0062", x"db6fe000", x"ec360000", x"f6bb6184", x"0aeb96e1", x"028686de", x"925e44c4"),
	(x"22860000", x"315e00ac", x"78b90000", x"93dc0000", x"8aff567c", x"959a9fea", x"f42553ad", x"715eb1d7", x"3ab70000", x"760d0074", x"c8330000", x"de2e0000", x"b8c0442c", x"6108e01e", x"c3667ecc", x"be0d07aa"),
	(x"a4ff0000", x"0e6700ae", x"9923e000", x"0b8a0000", x"1f9a3172", x"db125700", x"27f81ae9", x"67436b6e", x"0a000000", x"93dd0074", x"3cc76000", x"9cea0000", x"db787946", x"19b2747e", x"e2c9df26", x"0ea81f9e"),
	(x"12310000", x"d48e00ac", x"8c4d6000", x"d1180000", x"e9476b16", x"ed200b8a", x"d58af247", x"c1fba9e3", x"8c790000", x"ace40076", x"dd5d8000", x"04bc0000", x"4e1d1e48", x"573abc94", x"31149662", x"18b5c527"),
	(x"94480000", x"ebb700ae", x"6dd78000", x"494e0000", x"7c220c18", x"a3a8c360", x"0657bb03", x"d7e6735a", x"bcce0000", x"49340076", x"29a9e000", x"46780000", x"2da52322", x"2f8028f4", x"10bb3788", x"a810dd13"),
	(x"818c0000", x"2eab00d8", x"ff0e0000", x"173a0000", x"64283db5", x"ea4c0898", x"3844ea88", x"eeabae97", x"92230000", x"a9fc0050", x"816f0000", x"4b930000", x"0db45b58", x"1f5dd43d", x"a292b44b", x"49fc8c64"),
	(x"07f50000", x"119200da", x"1e94e000", x"8f6c0000", x"f14d5abb", x"a4c4c072", x"eb99a3cc", x"f8b6742e", x"a2940000", x"4c2c0050", x"759b6000", x"09570000", x"6e0c6632", x"67e7405d", x"833d15a1", x"f9599450"),
	(x"b13b0000", x"cb7b00d8", x"0bfa6000", x"55fe0000", x"079000df", x"92f69cf8", x"19eb4b62", x"5e0eb6a3", x"24ed0000", x"73150052", x"94018000", x"91010000", x"fb69013c", x"296f88b7", x"50e05ce5", x"ef444ee9"),
	(x"37420000", x"f44200da", x"ea608000", x"cda80000", x"92f567d1", x"dc7e5412", x"ca360226", x"48136c1a", x"145a0000", x"96c50052", x"60f5e000", x"d3c50000", x"98d13c56", x"51d51cd7", x"714ffd0f", x"5fe156dd"),
	(x"95950000", x"0d6100e4", x"afd10000", x"538c0000", x"7f445a05", x"d6bfa4ed", x"59a2fa38", x"35617517", x"71600000", x"93b20044", x"73a90000", x"e1dd0000", x"d6aa19fe", x"3a366a28", x"b0af051d", x"73b215b3"),
	(x"13ec0000", x"325800e6", x"4e4be000", x"cbda0000", x"ea213d0b", x"98376c07", x"8a7fb37c", x"237cafae", x"41d70000", x"76620044", x"875d6000", x"a3190000", x"b5122494", x"428cfe48", x"9100a4f7", x"c3170d87"),
	(x"a5220000", x"e8b100e4", x"5b256000", x"11480000", x"1cfc676f", x"ae05308d", x"780d5bd2", x"85c46d23", x"c7ae0000", x"495b0046", x"66c78000", x"3b4f0000", x"2077439a", x"0c0436a2", x"42ddedb3", x"d50ad73e"),
	(x"235b0000", x"d78800e6", x"babf8000", x"891e0000", x"89990061", x"e08df867", x"abd01296", x"93d9b79a", x"f7190000", x"ac8b0046", x"9233e000", x"798b0000", x"43cf7ef0", x"74bea2c2", x"63724c59", x"65afcf0a"),
	(x"62cf0000", x"14e500cc", x"0dc80000", x"bd740000", x"bf367f13", x"cf27b68d", x"2a795bde", x"d4e53740", x"65790000", x"b0780078", x"23760000", x"a56b0000", x"cdc67e4e", x"06c5c65d", x"d14915ad", x"a878ce33"),
	(x"e4b60000", x"2bdc00ce", x"ec52e000", x"25220000", x"2a53181d", x"81af7e67", x"f9a4129a", x"c2f8edf9", x"55ce0000", x"55a80078", x"d7826000", x"e7af0000", x"ae7e4324", x"7e7f523d", x"f0e6b447", x"18ddd607"),
	(x"52780000", x"f13500cc", x"f93c6000", x"ffb00000", x"dc8e4279", x"b79d22ed", x"0bd6fa34", x"64402f74", x"d3b70000", x"6a91007a", x"36188000", x"7ff90000", x"3b1b242a", x"30f79ad7", x"233bfd03", x"0ec00cbe"),
	(x"d4010000", x"ce0c00ce", x"18a68000", x"67e60000", x"49eb2577", x"f915ea07", x"d80bb370", x"725df5cd", x"e3000000", x"8f41007a", x"c2ece000", x"3d3d0000", x"58a31940", x"484d0eb7", x"02945ce9", x"be65148a"),
	(x"76d60000", x"372f00f0", x"5d170000", x"f9c20000", x"a45a18a3", x"f3d41af8", x"4b9f4b6e", x"0f2fecc0", x"863a0000", x"8a36006c", x"d1b00000", x"0f250000", x"16d83ce8", x"23ae7848", x"c374a4fb", x"923657e4"),
	(x"f0af0000", x"081600f2", x"bc8de000", x"61940000", x"313f7fad", x"bd5cd212", x"9842022a", x"19323679", x"b68d0000", x"6fe6006c", x"25446000", x"4de10000", x"75600182", x"5b14ec28", x"e2db0511", x"22934fd0"),
	(x"46610000", x"d2ff00f0", x"a9e36000", x"bb060000", x"c7e225c9", x"8b6e8e98", x"6a30ea84", x"bf8af4f4", x"30f40000", x"50df006e", x"c4de8000", x"d5b70000", x"e005668c", x"159c24c2", x"31064c55", x"348e9569"),
	(x"c0180000", x"edc600f2", x"48798000", x"23500000", x"528742c7", x"c5e64672", x"b9eda3c0", x"a9972e4d", x"00430000", x"b50f006e", x"302ae000", x"97730000", x"83bd5be6", x"6d26b0a2", x"10a9edbf", x"842b8d5d"),
	(x"c6730000", x"af8d000c", x"a4c10000", x"218d0000", x"23111587", x"7913512f", x"1d28ac88", x"378dd173", x"af220000", x"7b6c0090", x"67e20000", x"8da20000", x"c7841e29", x"b7b744f3", x"9ac484f4", x"8b6c72bd"),
	(x"400a0000", x"90b4000e", x"455be000", x"b9db0000", x"b6747289", x"379b99c5", x"cef5e5cc", x"21900bca", x"9f950000", x"9ebc0090", x"93166000", x"cf660000", x"a43c2343", x"cf0dd093", x"bb6b251e", x"3bc96a89"),
	(x"f6c40000", x"4a5d000c", x"50356000", x"63490000", x"40a928ed", x"01a9c54f", x"3c870d62", x"8728c947", x"19ec0000", x"a1850092", x"728c8000", x"57300000", x"3159444d", x"81851879", x"68b66c5a", x"2dd4b030"),
	(x"70bd0000", x"7564000e", x"b1af8000", x"fb1f0000", x"d5cc4fe3", x"4f210da5", x"ef5a4426", x"913513fe", x"295b0000", x"44550092", x"8678e000", x"15f40000", x"52e17927", x"f93f8c19", x"4919cdb0", x"9d71a804"),
	(x"d26a0000", x"8c470030", x"f41e0000", x"653b0000", x"387d7237", x"45e0fd5a", x"7ccebc38", x"ec470af3", x"4c610000", x"41220084", x"95240000", x"27ec0000", x"1c9a5c8f", x"92dcfae6", x"88f935a2", x"b122eb6a"),
	(x"54130000", x"b37e0032", x"1584e000", x"fd6d0000", x"ad181539", x"0b6835b0", x"af13f57c", x"fa5ad04a", x"7cd60000", x"a4f20084", x"61d06000", x"65280000", x"7f2261e5", x"ea666e86", x"a9569448", x"0187f35e"),
	(x"e2dd0000", x"69970030", x"00ea6000", x"27ff0000", x"5bc54f5d", x"3d5a693a", x"5d611dd2", x"5ce212c7", x"faaf0000", x"9bcb0086", x"804a8000", x"fd7e0000", x"ea4706eb", x"a4eea66c", x"7a8bdd0c", x"179a29e7"),
	(x"64a40000", x"56ae0032", x"e1708000", x"bfa90000", x"cea02853", x"73d2a1d0", x"8ebc5496", x"4affc87e", x"ca180000", x"7e1b0086", x"74bee000", x"bfba0000", x"89ff3b81", x"dc54320c", x"5b247ce6", x"a73f31d3"),
	(x"25300000", x"95c30018", x"56070000", x"8bc30000", x"f80f5721", x"5c78ef3a", x"0f151dde", x"0dc348a4", x"58780000", x"62e800b8", x"c5fb0000", x"635a0000", x"07f63b3f", x"ae2f5693", x"e91f2512", x"6ae830ea"),
	(x"a3490000", x"aafa001a", x"b79de000", x"13950000", x"6d6a302f", x"12f027d0", x"dcc8549a", x"1bde921d", x"68cf0000", x"873800b8", x"310f6000", x"219e0000", x"644e0655", x"d695c2f3", x"c8b084f8", x"da4d28de"),
	(x"15870000", x"70130018", x"a2f36000", x"c9070000", x"9bb76a4b", x"24c27b5a", x"2ebabc34", x"bd665090", x"eeb60000", x"b80100ba", x"d0958000", x"b9c80000", x"f12b615b", x"981d0a19", x"1b6dcdbc", x"cc50f267"),
	(x"93fe0000", x"4f2a001a", x"43698000", x"51510000", x"0ed20d45", x"6a4ab3b0", x"fd67f570", x"ab7b8a29", x"de010000", x"5dd100ba", x"2461e000", x"fb0c0000", x"92935c31", x"e0a79e79", x"3ac26c56", x"7cf5ea53"),
	(x"31290000", x"b6090024", x"06d80000", x"cf750000", x"e3633091", x"608b434f", x"6ef30d6e", x"d6099324", x"bb3b0000", x"58a600ac", x"373d0000", x"c9140000", x"dce87999", x"8b44e886", x"fb229444", x"50a6a93d"),
	(x"b7500000", x"89300026", x"e742e000", x"57230000", x"7606579f", x"2e038ba5", x"bd2e442a", x"c014499d", x"8b8c0000", x"bd7600ac", x"c3c96000", x"8bd00000", x"bf5044f3", x"f3fe7ce6", x"da8d35ae", x"e003b109"),
	(x"019e0000", x"53d90024", x"f22c6000", x"8db10000", x"80db0dfb", x"1831d72f", x"4f5cac84", x"66ac8b10", x"0df50000", x"824f00ae", x"22538000", x"13860000", x"2a3523fd", x"bd76b40c", x"09507cea", x"f61e6bb0"),
	(x"87e70000", x"6ce00026", x"13b68000", x"15e70000", x"15be6af5", x"56b91fc5", x"9c81e5c0", x"70b151a9", x"3d420000", x"679f00ae", x"d6a7e000", x"51420000", x"498d1e97", x"c5cc206c", x"28ffdd00", x"46bb7384"),
	(x"92230000", x"a9fc0050", x"816f0000", x"4b930000", x"0db45b58", x"1f5dd43d", x"a292b44b", x"49fc8c64", x"13af0000", x"87570088", x"7e610000", x"5ca90000", x"699c66ed", x"f511dca5", x"9ad65ec3", x"a75722f3"),
	(x"145a0000", x"96c50052", x"60f5e000", x"d3c50000", x"98d13c56", x"51d51cd7", x"714ffd0f", x"5fe156dd", x"23180000", x"62870088", x"8a956000", x"1e6d0000", x"0a245b87", x"8dab48c5", x"bb79ff29", x"17f23ac7"),
	(x"a2940000", x"4c2c0050", x"759b6000", x"09570000", x"6e0c6632", x"67e7405d", x"833d15a1", x"f9599450", x"a5610000", x"5dbe008a", x"6b0f8000", x"863b0000", x"9f413c89", x"c323802f", x"68a4b66d", x"01efe07e"),
	(x"24ed0000", x"73150052", x"94018000", x"91010000", x"fb69013c", x"296f88b7", x"50e05ce5", x"ef444ee9", x"95d60000", x"b86e008a", x"9ffbe000", x"c4ff0000", x"fcf901e3", x"bb99144f", x"490b1787", x"b14af84a"),
	(x"863a0000", x"8a36006c", x"d1b00000", x"0f250000", x"16d83ce8", x"23ae7848", x"c374a4fb", x"923657e4", x"f0ec0000", x"bd19009c", x"8ca70000", x"f6e70000", x"b282244b", x"d07a62b0", x"88ebef95", x"9d19bb24"),
	(x"00430000", x"b50f006e", x"302ae000", x"97730000", x"83bd5be6", x"6d26b0a2", x"10a9edbf", x"842b8d5d", x"c05b0000", x"58c9009c", x"78536000", x"b4230000", x"d13a1921", x"a8c0f6d0", x"a9444e7f", x"2dbca310"),
	(x"b68d0000", x"6fe6006c", x"25446000", x"4de10000", x"75600182", x"5b14ec28", x"e2db0511", x"22934fd0", x"46220000", x"67f0009e", x"99c98000", x"2c750000", x"445f7e2f", x"e6483e3a", x"7a99073b", x"3ba179a9"),
	(x"30f40000", x"50df006e", x"c4de8000", x"d5b70000", x"e005668c", x"159c24c2", x"31064c55", x"348e9569", x"76950000", x"8220009e", x"6d3de000", x"6eb10000", x"27e74345", x"9ef2aa5a", x"5b36a6d1", x"8b04619d"),
	(x"71600000", x"93b20044", x"73a90000", x"e1dd0000", x"d6aa19fe", x"3a366a28", x"b0af051d", x"73b215b3", x"e4f50000", x"9ed300a0", x"dc780000", x"b2510000", x"a9ee43fb", x"ec89cec5", x"e90dff25", x"46d360a4"),
	(x"f7190000", x"ac8b0046", x"9233e000", x"798b0000", x"43cf7ef0", x"74bea2c2", x"63724c59", x"65afcf0a", x"d4420000", x"7b0300a0", x"288c6000", x"f0950000", x"ca567e91", x"94335aa5", x"c8a25ecf", x"f6767890"),
	(x"41d70000", x"76620044", x"875d6000", x"a3190000", x"b5122494", x"428cfe48", x"9100a4f7", x"c3170d87", x"523b0000", x"443a00a2", x"c9168000", x"68c30000", x"5f33199f", x"dabb924f", x"1b7f178b", x"e06ba229"),
	(x"c7ae0000", x"495b0046", x"66c78000", x"3b4f0000", x"2077439a", x"0c0436a2", x"42ddedb3", x"d50ad73e", x"628c0000", x"a1ea00a2", x"3de2e000", x"2a070000", x"3c8b24f5", x"a201062f", x"3ad0b661", x"50ceba1d"),
	(x"65790000", x"b0780078", x"23760000", x"a56b0000", x"cdc67e4e", x"06c5c65d", x"d14915ad", x"a878ce33", x"07b60000", x"a49d00b4", x"2ebe0000", x"181f0000", x"72f0015d", x"c9e270d0", x"fb304e73", x"7c9df973"),
	(x"e3000000", x"8f41007a", x"c2ece000", x"3d3d0000", x"58a31940", x"484d0eb7", x"02945ce9", x"be65148a", x"37010000", x"414d00b4", x"da4a6000", x"5adb0000", x"11483c37", x"b158e4b0", x"da9fef99", x"cc38e147"),
	(x"55ce0000", x"55a80078", x"d7826000", x"e7af0000", x"ae7e4324", x"7e7f523d", x"f0e6b447", x"18ddd607", x"b1780000", x"7e7400b6", x"3bd08000", x"c28d0000", x"842d5b39", x"ffd02c5a", x"0942a6dd", x"da253bfe"),
	(x"d3b70000", x"6a91007a", x"36188000", x"7ff90000", x"3b1b242a", x"30f79ad7", x"233bfd03", x"0ec00cbe", x"81cf0000", x"9ba400b6", x"cf24e000", x"80490000", x"e7956653", x"876ab83a", x"28ed0737", x"6a8023ca"),
	(x"7afe0000", x"53b60014", x"bd420000", x"f0860000", x"8d096d43", x"3bb5c979", x"1d3a76bf", x"1bb6813d", x"47ff0000", x"812600d4", x"5bcf0000", x"36b70000", x"47392832", x"935f59b7", x"256c4600", x"d9267fe4"),
	(x"fc870000", x"6c8f0016", x"5cd8e000", x"68d00000", x"186c0a4d", x"753d0193", x"cee73ffb", x"0dab5b84", x"77480000", x"64f600d4", x"af3b6000", x"74730000", x"24811558", x"ebe5cdd7", x"04c3e7ea", x"698367d0"),
	(x"4a490000", x"b6660014", x"49b66000", x"b2420000", x"eeb15029", x"430f5d19", x"3c95d755", x"ab139909", x"f1310000", x"5bcf00d6", x"4ea18000", x"ec250000", x"b1e47256", x"a56d053d", x"d71eaeae", x"7f9ebd69"),
	(x"cc300000", x"895f0016", x"a82c8000", x"2a140000", x"7bd43727", x"0d8795f3", x"ef489e11", x"bd0e43b0", x"c1860000", x"be1f00d6", x"ba55e000", x"aee10000", x"d25c4f3c", x"ddd7915d", x"f6b10f44", x"cf3ba55d"),
	(x"6ee70000", x"707c0028", x"ed9d0000", x"b4300000", x"96650af3", x"0746650c", x"7cdc660f", x"c07c5abd", x"a4bc0000", x"bb6800c0", x"a9090000", x"9cf90000", x"9c276a94", x"b634e7a2", x"3751f756", x"e368e633"),
	(x"e89e0000", x"4f45002a", x"0c07e000", x"2c660000", x"03006dfd", x"49ceade6", x"af012f4b", x"d6618004", x"940b0000", x"5eb800c0", x"5dfd6000", x"de3d0000", x"ff9f57fe", x"ce8e73c2", x"16fe56bc", x"53cdfe07"),
	(x"5e500000", x"95ac0028", x"19696000", x"f6f40000", x"f5dd3799", x"7ffcf16c", x"5d73c7e5", x"70d94289", x"12720000", x"618100c2", x"bc678000", x"466b0000", x"6afa30f0", x"8006bb28", x"c5231ff8", x"45d024be"),
	(x"d8290000", x"aa95002a", x"f8f38000", x"6ea20000", x"60b85097", x"31743986", x"8eae8ea1", x"66c49830", x"22c50000", x"845100c2", x"4893e000", x"04af0000", x"09420d9a", x"f8bc2f48", x"e48cbe12", x"f5753c8a"),
	(x"99bd0000", x"69f80000", x"4f840000", x"5ac80000", x"56172fe5", x"1ede776c", x"0f07c7e9", x"21f818ea", x"b0a50000", x"98a200fc", x"f9d60000", x"d84f0000", x"874b0d24", x"8ac74bd7", x"56b7e7e6", x"38a23db3"),
	(x"1fc40000", x"56c10002", x"ae1ee000", x"c29e0000", x"c37248eb", x"5056bf86", x"dcda8ead", x"37e5c253", x"80120000", x"7d7200fc", x"0d226000", x"9a8b0000", x"e4f3304e", x"f27ddfb7", x"7718460c", x"88072587"),
	(x"a90a0000", x"8c280000", x"bb706000", x"180c0000", x"35af128f", x"6664e30c", x"2ea86603", x"915d00de", x"066b0000", x"424b00fe", x"ecb88000", x"02dd0000", x"71965740", x"bcf5175d", x"a4c50f48", x"9e1aff3e"),
	(x"2f730000", x"b3110002", x"5aea8000", x"805a0000", x"a0ca7581", x"28ec2be6", x"fd752f47", x"8740da67", x"36dc0000", x"a79b00fe", x"184ce000", x"40190000", x"122e6a2a", x"c44f833d", x"856aaea2", x"2ebfe70a"),
	(x"8da40000", x"4a32003c", x"1f5b0000", x"1e7e0000", x"4d7b4855", x"222ddb19", x"6ee1d759", x"fa32c36a", x"53e60000", x"a2ec00e8", x"0b100000", x"72010000", x"5c554f82", x"afacf5c2", x"448a56b0", x"02eca464"),
	(x"0bdd0000", x"750b003e", x"fec1e000", x"86280000", x"d81e2f5b", x"6ca513f3", x"bd3c9e1d", x"ec2f19d3", x"63510000", x"473c00e8", x"ffe46000", x"30c50000", x"3fed72e8", x"d71661a2", x"6525f75a", x"b249bc50"),
	(x"bd130000", x"afe2003c", x"ebaf6000", x"5cba0000", x"2ec3753f", x"5a974f79", x"4f4e76b3", x"4a97db5e", x"e5280000", x"780500ea", x"1e7e8000", x"a8930000", x"aa8815e6", x"999ea948", x"b6f8be1e", x"a45466e9"),
	(x"3b6a0000", x"90db003e", x"0a358000", x"c4ec0000", x"bba61231", x"141f8793", x"9c933ff7", x"5c8a01e7", x"d59f0000", x"9dd500ea", x"ea8ae000", x"ea570000", x"c930288c", x"e1243d28", x"97571ff4", x"14f17edd"),
	(x"2eae0000", x"55c70048", x"98ec0000", x"9a980000", x"a3ac239c", x"5dfb4c6b", x"a2806e7c", x"65c7dc2a", x"fb720000", x"7d1d00cc", x"424c0000", x"e7bc0000", x"e92150f6", x"d1f9c1e1", x"257e9c37", x"f51d2faa"),
	(x"a8d70000", x"6afe004a", x"7976e000", x"02ce0000", x"36c94492", x"13738481", x"715d2738", x"73da0693", x"cbc50000", x"98cd00cc", x"b6b86000", x"a5780000", x"8a996d9c", x"a9435581", x"04d13ddd", x"45b8379e"),
	(x"1e190000", x"b0170048", x"6c186000", x"d85c0000", x"c0141ef6", x"2541d80b", x"832fcf96", x"d562c41e", x"4dbc0000", x"a7f400ce", x"57228000", x"3d2e0000", x"1ffc0a92", x"e7cb9d6b", x"d70c7499", x"53a5ed27"),
	(x"98600000", x"8f2e004a", x"8d828000", x"400a0000", x"557179f8", x"6bc910e1", x"50f286d2", x"c37f1ea7", x"7d0b0000", x"422400ce", x"a3d6e000", x"7fea0000", x"7c4437f8", x"9f71090b", x"f6a3d573", x"e300f513"),
	(x"3ab70000", x"760d0074", x"c8330000", x"de2e0000", x"b8c0442c", x"6108e01e", x"c3667ecc", x"be0d07aa", x"18310000", x"475300d8", x"b08a0000", x"4df20000", x"323f1250", x"f4927ff4", x"37432d61", x"cf53b67d"),
	(x"bcce0000", x"49340076", x"29a9e000", x"46780000", x"2da52322", x"2f8028f4", x"10bb3788", x"a810dd13", x"28860000", x"a28300d8", x"447e6000", x"0f360000", x"51872f3a", x"8c28eb94", x"16ec8c8b", x"7ff6ae49"),
	(x"0a000000", x"93dd0074", x"3cc76000", x"9cea0000", x"db787946", x"19b2747e", x"e2c9df26", x"0ea81f9e", x"aeff0000", x"9dba00da", x"a5e48000", x"97600000", x"c4e24834", x"c2a0237e", x"c531c5cf", x"69eb74f0"),
	(x"8c790000", x"ace40076", x"dd5d8000", x"04bc0000", x"4e1d1e48", x"573abc94", x"31149662", x"18b5c527", x"9e480000", x"786a00da", x"5110e000", x"d5a40000", x"a75a755e", x"ba1ab71e", x"e49e6425", x"d94e6cc4"),
	(x"cded0000", x"6f89005c", x"6a2a0000", x"30d60000", x"78b2613a", x"7890f27e", x"b0bddf2a", x"5f8945fd", x"0c280000", x"649900e4", x"e0550000", x"09440000", x"295375e0", x"c861d381", x"56a53dd1", x"14996dfd"),
	(x"4b940000", x"50b0005e", x"8bb0e000", x"a8800000", x"edd70634", x"36183a94", x"6360966e", x"49949f44", x"3c9f0000", x"814900e4", x"14a16000", x"4b800000", x"4aeb488a", x"b0db47e1", x"770a9c3b", x"a43c75c9"),
	(x"fd5a0000", x"8a59005c", x"9ede6000", x"72120000", x"1b0a5c50", x"002a661e", x"91127ec0", x"ef2c5dc9", x"bae60000", x"be7000e6", x"f53b8000", x"d3d60000", x"df8e2f84", x"fe538f0b", x"a4d7d57f", x"b221af70"),
	(x"7b230000", x"b560005e", x"7f448000", x"ea440000", x"8e6f3b5e", x"4ea2aef4", x"42cf3784", x"f9318770", x"8a510000", x"5ba000e6", x"01cfe000", x"91120000", x"bc3612ee", x"86e91b6b", x"85787495", x"0284b744"),
	(x"d9f40000", x"4c430060", x"3af50000", x"74600000", x"63de068a", x"44635e0b", x"d15bcf9a", x"84439e7d", x"ef6b0000", x"5ed700f0", x"12930000", x"a30a0000", x"f24d3746", x"ed0a6d94", x"44988c87", x"2ed7f42a"),
	(x"5f8d0000", x"737a0062", x"db6fe000", x"ec360000", x"f6bb6184", x"0aeb96e1", x"028686de", x"925e44c4", x"dfdc0000", x"bb0700f0", x"e6676000", x"e1ce0000", x"91f50a2c", x"95b0f9f4", x"65372d6d", x"9e72ec1e"),
	(x"e9430000", x"a9930060", x"ce016000", x"36a40000", x"00663be0", x"3cd9ca6b", x"f0f46e70", x"34e68649", x"59a50000", x"843e00f2", x"07fd8000", x"79980000", x"04906d22", x"db38311e", x"b6ea6429", x"886f36a7"),
	(x"6f3a0000", x"96aa0062", x"2f9b8000", x"aef20000", x"95035cee", x"72510281", x"23292734", x"22fb5cf0", x"69120000", x"61ee00f2", x"f309e000", x"3b5c0000", x"67285048", x"a382a57e", x"9745c5c3", x"38ca2e93"),
	(x"af220000", x"7b6c0090", x"67e20000", x"8da20000", x"c7841e29", x"b7b744f3", x"9ac484f4", x"8b6c72bd", x"69510000", x"d4e1009c", x"c3230000", x"ac2f0000", x"e4950bae", x"cea415dc", x"87ec287c", x"bce1a3ce"),
	(x"295b0000", x"44550092", x"8678e000", x"15f40000", x"52e17927", x"f93f8c19", x"4919cdb0", x"9d71a804", x"59e60000", x"3131009c", x"37d76000", x"eeeb0000", x"872d36c4", x"b61e81bc", x"a6438996", x"0c44bbfa"),
	(x"9f950000", x"9ebc0090", x"93166000", x"cf660000", x"a43c2343", x"cf0dd093", x"bb6b251e", x"3bc96a89", x"df9f0000", x"0e08009e", x"d64d8000", x"76bd0000", x"124851ca", x"f8964956", x"759ec0d2", x"1a596143"),
	(x"19ec0000", x"a1850092", x"728c8000", x"57300000", x"3159444d", x"81851879", x"68b66c5a", x"2dd4b030", x"ef280000", x"ebd8009e", x"22b9e000", x"34790000", x"71f06ca0", x"802cdd36", x"54316138", x"aafc7977"),
	(x"bb3b0000", x"58a600ac", x"373d0000", x"c9140000", x"dce87999", x"8b44e886", x"fb229444", x"50a6a93d", x"8a120000", x"eeaf0088", x"31e50000", x"06610000", x"3f8b4908", x"ebcfabc9", x"95d1992a", x"86af3a19"),
	(x"3d420000", x"679f00ae", x"d6a7e000", x"51420000", x"498d1e97", x"c5cc206c", x"28ffdd00", x"46bb7384", x"baa50000", x"0b7f0088", x"c5116000", x"44a50000", x"5c337462", x"93753fa9", x"b47e38c0", x"360a222d"),
	(x"8b8c0000", x"bd7600ac", x"c3c96000", x"8bd00000", x"bf5044f3", x"f3fe7ce6", x"da8d35ae", x"e003b109", x"3cdc0000", x"3446008a", x"248b8000", x"dcf30000", x"c956136c", x"ddfdf743", x"67a37184", x"2017f894"),
	(x"0df50000", x"824f00ae", x"22538000", x"13860000", x"2a3523fd", x"bd76b40c", x"09507cea", x"f61e6bb0", x"0c6b0000", x"d196008a", x"d07fe000", x"9e370000", x"aaee2e06", x"a5476323", x"460cd06e", x"90b2e0a0"),
	(x"4c610000", x"41220084", x"95240000", x"27ec0000", x"1c9a5c8f", x"92dcfae6", x"88f935a2", x"b122eb6a", x"9e0b0000", x"cd6500b4", x"613a0000", x"42d70000", x"24e72eb8", x"d73c07bc", x"f437899a", x"5d65e199"),
	(x"ca180000", x"7e1b0086", x"74bee000", x"bfba0000", x"89ff3b81", x"dc54320c", x"5b247ce6", x"a73f31d3", x"aebc0000", x"28b500b4", x"95ce6000", x"00130000", x"475f13d2", x"af8693dc", x"d5982870", x"edc0f9ad"),
	(x"7cd60000", x"a4f20084", x"61d06000", x"65280000", x"7f2261e5", x"ea666e86", x"a9569448", x"0187f35e", x"28c50000", x"178c00b6", x"74548000", x"98450000", x"d23a74dc", x"e10e5b36", x"06456134", x"fbdd2314"),
	(x"faaf0000", x"9bcb0086", x"804a8000", x"fd7e0000", x"ea4706eb", x"a4eea66c", x"7a8bdd0c", x"179a29e7", x"18720000", x"f25c00b6", x"80a0e000", x"da810000", x"b18249b6", x"99b4cf56", x"27eac0de", x"4b783b20"),
	(x"58780000", x"62e800b8", x"c5fb0000", x"635a0000", x"07f63b3f", x"ae2f5693", x"e91f2512", x"6ae830ea", x"7d480000", x"f72b00a0", x"93fc0000", x"e8990000", x"fff96c1e", x"f257b9a9", x"e60a38cc", x"672b784e"),
	(x"de010000", x"5dd100ba", x"2461e000", x"fb0c0000", x"92935c31", x"e0a79e79", x"3ac26c56", x"7cf5ea53", x"4dff0000", x"12fb00a0", x"67086000", x"aa5d0000", x"9c415174", x"8aed2dc9", x"c7a59926", x"d78e607a"),
	(x"68cf0000", x"873800b8", x"310f6000", x"219e0000", x"644e0655", x"d695c2f3", x"c8b084f8", x"da4d28de", x"cb860000", x"2dc200a2", x"86928000", x"320b0000", x"0924367a", x"c465e523", x"1478d062", x"c193bac3"),
	(x"eeb60000", x"b80100ba", x"d0958000", x"b9c80000", x"f12b615b", x"981d0a19", x"1b6dcdbc", x"cc50f267", x"fb310000", x"c81200a2", x"7266e000", x"70cf0000", x"6a9c0b10", x"bcdf7143", x"35d77188", x"7136a2f7"),
	(x"fb720000", x"7d1d00cc", x"424c0000", x"e7bc0000", x"e92150f6", x"d1f9c1e1", x"257e9c37", x"f51d2faa", x"d5dc0000", x"28da0084", x"daa00000", x"7d240000", x"4a8d736a", x"8c028d8a", x"87fef24b", x"90daf380"),
	(x"7d0b0000", x"422400ce", x"a3d6e000", x"7fea0000", x"7c4437f8", x"9f71090b", x"f6a3d573", x"e300f513", x"e56b0000", x"cd0a0084", x"2e546000", x"3fe00000", x"29354e00", x"f4b819ea", x"a65153a1", x"207febb4"),
	(x"cbc50000", x"98cd00cc", x"b6b86000", x"a5780000", x"8a996d9c", x"a9435581", x"04d13ddd", x"45b8379e", x"63120000", x"f2330086", x"cfce8000", x"a7b60000", x"bc50290e", x"ba30d100", x"758c1ae5", x"3662310d"),
	(x"4dbc0000", x"a7f400ce", x"57228000", x"3d2e0000", x"1ffc0a92", x"e7cb9d6b", x"d70c7499", x"53a5ed27", x"53a50000", x"17e30086", x"3b3ae000", x"e5720000", x"dfe81464", x"c28a4560", x"5423bb0f", x"86c72939"),
	(x"ef6b0000", x"5ed700f0", x"12930000", x"a30a0000", x"f24d3746", x"ed0a6d94", x"44988c87", x"2ed7f42a", x"369f0000", x"12940090", x"28660000", x"d76a0000", x"919331cc", x"a969339f", x"95c3431d", x"aa946a57"),
	(x"69120000", x"61ee00f2", x"f309e000", x"3b5c0000", x"67285048", x"a382a57e", x"9745c5c3", x"38ca2e93", x"06280000", x"f7440090", x"dc926000", x"95ae0000", x"f22b0ca6", x"d1d3a7ff", x"b46ce2f7", x"1a317263"),
	(x"dfdc0000", x"bb0700f0", x"e6676000", x"e1ce0000", x"91f50a2c", x"95b0f9f4", x"65372d6d", x"9e72ec1e", x"80510000", x"c87d0092", x"3d088000", x"0df80000", x"674e6ba8", x"9f5b6f15", x"67b1abb3", x"0c2ca8da"),
	(x"59a50000", x"843e00f2", x"07fd8000", x"79980000", x"04906d22", x"db38311e", x"b6ea6429", x"886f36a7", x"b0e60000", x"2dad0092", x"c9fce000", x"4f3c0000", x"04f656c2", x"e7e1fb75", x"461e0a59", x"bc89b0ee"),
	(x"18310000", x"475300d8", x"b08a0000", x"4df20000", x"323f1250", x"f4927ff4", x"37432d61", x"cf53b67d", x"22860000", x"315e00ac", x"78b90000", x"93dc0000", x"8aff567c", x"959a9fea", x"f42553ad", x"715eb1d7"),
	(x"9e480000", x"786a00da", x"5110e000", x"d5a40000", x"a75a755e", x"ba1ab71e", x"e49e6425", x"d94e6cc4", x"12310000", x"d48e00ac", x"8c4d6000", x"d1180000", x"e9476b16", x"ed200b8a", x"d58af247", x"c1fba9e3"),
	(x"28860000", x"a28300d8", x"447e6000", x"0f360000", x"51872f3a", x"8c28eb94", x"16ec8c8b", x"7ff6ae49", x"94480000", x"ebb700ae", x"6dd78000", x"494e0000", x"7c220c18", x"a3a8c360", x"0657bb03", x"d7e6735a"),
	(x"aeff0000", x"9dba00da", x"a5e48000", x"97600000", x"c4e24834", x"c2a0237e", x"c531c5cf", x"69eb74f0", x"a4ff0000", x"0e6700ae", x"9923e000", x"0b8a0000", x"1f9a3172", x"db125700", x"27f81ae9", x"67436b6e"),
	(x"0c280000", x"649900e4", x"e0550000", x"09440000", x"295375e0", x"c861d381", x"56a53dd1", x"14996dfd", x"c1c50000", x"0b1000b8", x"8a7f0000", x"39920000", x"51e114da", x"b0f121ff", x"e618e2fb", x"4b102800"),
	(x"8a510000", x"5ba000e6", x"01cfe000", x"91120000", x"bc3612ee", x"86e91b6b", x"85787495", x"0284b744", x"f1720000", x"eec000b8", x"7e8b6000", x"7b560000", x"325929b0", x"c84bb59f", x"c7b74311", x"fbb53034"),
	(x"3c9f0000", x"814900e4", x"14a16000", x"4b800000", x"4aeb488a", x"b0db47e1", x"770a9c3b", x"a43c75c9", x"770b0000", x"d1f900ba", x"9f118000", x"e3000000", x"a73c4ebe", x"86c37d75", x"146a0a55", x"eda8ea8d"),
	(x"bae60000", x"be7000e6", x"f53b8000", x"d3d60000", x"df8e2f84", x"fe538f0b", x"a4d7d57f", x"b221af70", x"47bc0000", x"342900ba", x"6be5e000", x"a1c40000", x"c48473d4", x"fe79e915", x"35c5abbf", x"5d0df2b9"),
	(x"13af0000", x"87570088", x"7e610000", x"5ca90000", x"699c66ed", x"f511dca5", x"9ad65ec3", x"a75722f3", x"818c0000", x"2eab00d8", x"ff0e0000", x"173a0000", x"64283db5", x"ea4c0898", x"3844ea88", x"eeabae97"),
	(x"95d60000", x"b86e008a", x"9ffbe000", x"c4ff0000", x"fcf901e3", x"bb99144f", x"490b1787", x"b14af84a", x"b13b0000", x"cb7b00d8", x"0bfa6000", x"55fe0000", x"079000df", x"92f69cf8", x"19eb4b62", x"5e0eb6a3"),
	(x"23180000", x"62870088", x"8a956000", x"1e6d0000", x"0a245b87", x"8dab48c5", x"bb79ff29", x"17f23ac7", x"37420000", x"f44200da", x"ea608000", x"cda80000", x"92f567d1", x"dc7e5412", x"ca360226", x"48136c1a"),
	(x"a5610000", x"5dbe008a", x"6b0f8000", x"863b0000", x"9f413c89", x"c323802f", x"68a4b66d", x"01efe07e", x"07f50000", x"119200da", x"1e94e000", x"8f6c0000", x"f14d5abb", x"a4c4c072", x"eb99a3cc", x"f8b6742e"),
	(x"07b60000", x"a49d00b4", x"2ebe0000", x"181f0000", x"72f0015d", x"c9e270d0", x"fb304e73", x"7c9df973", x"62cf0000", x"14e500cc", x"0dc80000", x"bd740000", x"bf367f13", x"cf27b68d", x"2a795bde", x"d4e53740"),
	(x"81cf0000", x"9ba400b6", x"cf24e000", x"80490000", x"e7956653", x"876ab83a", x"28ed0737", x"6a8023ca", x"52780000", x"f13500cc", x"f93c6000", x"ffb00000", x"dc8e4279", x"b79d22ed", x"0bd6fa34", x"64402f74"),
	(x"37010000", x"414d00b4", x"da4a6000", x"5adb0000", x"11483c37", x"b158e4b0", x"da9fef99", x"cc38e147", x"d4010000", x"ce0c00ce", x"18a68000", x"67e60000", x"49eb2577", x"f915ea07", x"d80bb370", x"725df5cd"),
	(x"b1780000", x"7e7400b6", x"3bd08000", x"c28d0000", x"842d5b39", x"ffd02c5a", x"0942a6dd", x"da253bfe", x"e4b60000", x"2bdc00ce", x"ec52e000", x"25220000", x"2a53181d", x"81af7e67", x"f9a4129a", x"c2f8edf9"),
	(x"f0ec0000", x"bd19009c", x"8ca70000", x"f6e70000", x"b282244b", x"d07a62b0", x"88ebef95", x"9d19bb24", x"76d60000", x"372f00f0", x"5d170000", x"f9c20000", x"a45a18a3", x"f3d41af8", x"4b9f4b6e", x"0f2fecc0"),
	(x"76950000", x"8220009e", x"6d3de000", x"6eb10000", x"27e74345", x"9ef2aa5a", x"5b36a6d1", x"8b04619d", x"46610000", x"d2ff00f0", x"a9e36000", x"bb060000", x"c7e225c9", x"8b6e8e98", x"6a30ea84", x"bf8af4f4"),
	(x"c05b0000", x"58c9009c", x"78536000", x"b4230000", x"d13a1921", x"a8c0f6d0", x"a9444e7f", x"2dbca310", x"c0180000", x"edc600f2", x"48798000", x"23500000", x"528742c7", x"c5e64672", x"b9eda3c0", x"a9972e4d"),
	(x"46220000", x"67f0009e", x"99c98000", x"2c750000", x"445f7e2f", x"e6483e3a", x"7a99073b", x"3ba179a9", x"f0af0000", x"081600f2", x"bc8de000", x"61940000", x"313f7fad", x"bd5cd212", x"9842022a", x"19323679"),
	(x"e4f50000", x"9ed300a0", x"dc780000", x"b2510000", x"a9ee43fb", x"ec89cec5", x"e90dff25", x"46d360a4", x"95950000", x"0d6100e4", x"afd10000", x"538c0000", x"7f445a05", x"d6bfa4ed", x"59a2fa38", x"35617517"),
	(x"628c0000", x"a1ea00a2", x"3de2e000", x"2a070000", x"3c8b24f5", x"a201062f", x"3ad0b661", x"50ceba1d", x"a5220000", x"e8b100e4", x"5b256000", x"11480000", x"1cfc676f", x"ae05308d", x"780d5bd2", x"85c46d23"),
	(x"d4420000", x"7b0300a0", x"288c6000", x"f0950000", x"ca567e91", x"94335aa5", x"c8a25ecf", x"f6767890", x"235b0000", x"d78800e6", x"babf8000", x"891e0000", x"89990061", x"e08df867", x"abd01296", x"93d9b79a"),
	(x"523b0000", x"443a00a2", x"c9168000", x"68c30000", x"5f33199f", x"dabb924f", x"1b7f178b", x"e06ba229", x"13ec0000", x"325800e6", x"4e4be000", x"cbda0000", x"ea213d0b", x"98376c07", x"8a7fb37c", x"237cafae"),
	(x"47ff0000", x"812600d4", x"5bcf0000", x"36b70000", x"47392832", x"935f59b7", x"256c4600", x"d9267fe4", x"3d010000", x"d29000c0", x"e68d0000", x"c6310000", x"ca304571", x"a8ea90ce", x"385630bf", x"c290fed9"),
	(x"c1860000", x"be1f00d6", x"ba55e000", x"aee10000", x"d25c4f3c", x"ddd7915d", x"f6b10f44", x"cf3ba55d", x"0db60000", x"374000c0", x"12796000", x"84f50000", x"a988781b", x"d05004ae", x"19f99155", x"7235e6ed"),
	(x"77480000", x"64f600d4", x"af3b6000", x"74730000", x"24811558", x"ebe5cdd7", x"04c3e7ea", x"698367d0", x"8bcf0000", x"087900c2", x"f3e38000", x"1ca30000", x"3ced1f15", x"9ed8cc44", x"ca24d811", x"64283c54"),
	(x"f1310000", x"5bcf00d6", x"4ea18000", x"ec250000", x"b1e47256", x"a56d053d", x"d71eaeae", x"7f9ebd69", x"bb780000", x"eda900c2", x"0717e000", x"5e670000", x"5f55227f", x"e6625824", x"eb8b79fb", x"d48d2460"),
	(x"53e60000", x"a2ec00e8", x"0b100000", x"72010000", x"5c554f82", x"afacf5c2", x"448a56b0", x"02eca464", x"de420000", x"e8de00d4", x"144b0000", x"6c7f0000", x"112e07d7", x"8d812edb", x"2a6b81e9", x"f8de670e"),
	(x"d59f0000", x"9dd500ea", x"ea8ae000", x"ea570000", x"c930288c", x"e1243d28", x"97571ff4", x"14f17edd", x"eef50000", x"0d0e00d4", x"e0bf6000", x"2ebb0000", x"72963abd", x"f53bbabb", x"0bc42003", x"487b7f3a"),
	(x"63510000", x"473c00e8", x"ffe46000", x"30c50000", x"3fed72e8", x"d71661a2", x"6525f75a", x"b249bc50", x"688c0000", x"323700d6", x"01258000", x"b6ed0000", x"e7f35db3", x"bbb37251", x"d8196947", x"5e66a583"),
	(x"e5280000", x"780500ea", x"1e7e8000", x"a8930000", x"aa8815e6", x"999ea948", x"b6f8be1e", x"a45466e9", x"583b0000", x"d7e700d6", x"f5d1e000", x"f4290000", x"844b60d9", x"c309e631", x"f9b6c8ad", x"eec3bdb7"),
	(x"a4bc0000", x"bb6800c0", x"a9090000", x"9cf90000", x"9c276a94", x"b634e7a2", x"3751f756", x"e368e633", x"ca5b0000", x"cb1400e8", x"44940000", x"28c90000", x"0a426067", x"b17282ae", x"4b8d9159", x"2314bc8e"),
	(x"22c50000", x"845100c2", x"4893e000", x"04af0000", x"09420d9a", x"f8bc2f48", x"e48cbe12", x"f5753c8a", x"faec0000", x"2ec400e8", x"b0606000", x"6a0d0000", x"69fa5d0d", x"c9c816ce", x"6a2230b3", x"93b1a4ba"),
	(x"940b0000", x"5eb800c0", x"5dfd6000", x"de3d0000", x"ff9f57fe", x"ce8e73c2", x"16fe56bc", x"53cdfe07", x"7c950000", x"11fd00ea", x"51fa8000", x"f25b0000", x"fc9f3a03", x"8740de24", x"b9ff79f7", x"85ac7e03"),
	(x"12720000", x"618100c2", x"bc678000", x"466b0000", x"6afa30f0", x"8006bb28", x"c5231ff8", x"45d024be", x"4c220000", x"f42d00ea", x"a50ee000", x"b09f0000", x"9f270769", x"fffa4a44", x"9850d81d", x"35096637"),
	(x"b0a50000", x"98a200fc", x"f9d60000", x"d84f0000", x"874b0d24", x"8ac74bd7", x"56b7e7e6", x"38a23db3", x"29180000", x"f15a00fc", x"b6520000", x"82870000", x"d15c22c1", x"94193cbb", x"59b0200f", x"195a2559"),
	(x"36dc0000", x"a79b00fe", x"184ce000", x"40190000", x"122e6a2a", x"c44f833d", x"856aaea2", x"2ebfe70a", x"19af0000", x"148a00fc", x"42a66000", x"c0430000", x"b2e41fab", x"eca3a8db", x"781f81e5", x"a9ff3d6d"),
	(x"80120000", x"7d7200fc", x"0d226000", x"9a8b0000", x"e4f3304e", x"f27ddfb7", x"7718460c", x"88072587", x"9fd60000", x"2bb300fe", x"a33c8000", x"58150000", x"278178a5", x"a22b6031", x"abc2c8a1", x"bfe2e7d4"),
	(x"066b0000", x"424b00fe", x"ecb88000", x"02dd0000", x"71965740", x"bcf5175d", x"a4c50f48", x"9e1aff3e", x"af610000", x"ce6300fe", x"57c8e000", x"1ad10000", x"443945cf", x"da91f451", x"8a6d694b", x"0f47ffe0")
    ),(
	(x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000"),
	(x"cc140000", x"a5630000", x"5ab90780", x"3b500000", x"4bd013ff", x"879b3418", x"694348c1", x"ca5a87fe", x"819e0000", x"ec570000", x"66320280", x"95f30000", x"5da92802", x"48f43cbc", x"e65aa22d", x"8e67b7fa"),
	(x"819e0000", x"ec570000", x"66320280", x"95f30000", x"5da92802", x"48f43cbc", x"e65aa22d", x"8e67b7fa", x"4d8a0000", x"49340000", x"3c8b0500", x"aea30000", x"16793bfd", x"cf6f08a4", x"8f19eaec", x"443d3004"),
	(x"4d8a0000", x"49340000", x"3c8b0500", x"aea30000", x"16793bfd", x"cf6f08a4", x"8f19eaec", x"443d3004", x"cc140000", x"a5630000", x"5ab90780", x"3b500000", x"4bd013ff", x"879b3418", x"694348c1", x"ca5a87fe"),
	(x"78230000", x"12fc0000", x"a93a0b80", x"90a50000", x"713e2879", x"7ee98924", x"f08ca062", x"636f8bab", x"02af0000", x"b7280000", x"ba1c0300", x"56980000", x"ba8d45d3", x"8048c667", x"a95c149a", x"f4f6ea7b"),
	(x"b4370000", x"b79f0000", x"f3830c00", x"abf50000", x"3aee3b86", x"f972bd3c", x"99cfe8a3", x"a9350c55", x"83310000", x"5b7f0000", x"dc2e0180", x"c36b0000", x"e7246dd1", x"c8bcfadb", x"4f06b6b7", x"7a915d81"),
	(x"f9bd0000", x"feab0000", x"cf080900", x"05560000", x"2c97007b", x"361db598", x"16d6024f", x"ed083c51", x"4f250000", x"fe1c0000", x"86970600", x"f83b0000", x"acf47e2e", x"4f27cec3", x"2645fe76", x"b0cbda7f"),
	(x"35a90000", x"5bc80000", x"95b10e80", x"3e060000", x"67471384", x"b1868180", x"7f954a8e", x"2752bbaf", x"cebb0000", x"124b0000", x"e0a50480", x"6dc80000", x"f15d562c", x"07d3f27f", x"c01f5c5b", x"3eac6d85"),
	(x"02af0000", x"b7280000", x"ba1c0300", x"56980000", x"ba8d45d3", x"8048c667", x"a95c149a", x"f4f6ea7b", x"7a8c0000", x"a5d40000", x"13260880", x"c63d0000", x"cbb36daa", x"fea14f43", x"59d0b4f8", x"979961d0"),
	(x"cebb0000", x"124b0000", x"e0a50480", x"6dc80000", x"f15d562c", x"07d3f27f", x"c01f5c5b", x"3eac6d85", x"fb120000", x"49830000", x"75140a00", x"53ce0000", x"961a45a8", x"b65573ff", x"bf8a16d5", x"19fed62a"),
	(x"83310000", x"5b7f0000", x"dc2e0180", x"c36b0000", x"e7246dd1", x"c8bcfadb", x"4f06b6b7", x"7a915d81", x"37060000", x"ece00000", x"2fad0d80", x"689e0000", x"ddca5657", x"31ce47e7", x"d6c95e14", x"d3a451d4"),
	(x"4f250000", x"fe1c0000", x"86970600", x"f83b0000", x"acf47e2e", x"4f27cec3", x"2645fe76", x"b0cbda7f", x"b6980000", x"00b70000", x"499f0f00", x"fd6d0000", x"80637e55", x"793a7b5b", x"3093fc39", x"5dc3e62e"),
	(x"7a8c0000", x"a5d40000", x"13260880", x"c63d0000", x"cbb36daa", x"fea14f43", x"59d0b4f8", x"979961d0", x"78230000", x"12fc0000", x"a93a0b80", x"90a50000", x"713e2879", x"7ee98924", x"f08ca062", x"636f8bab"),
	(x"b6980000", x"00b70000", x"499f0f00", x"fd6d0000", x"80637e55", x"793a7b5b", x"3093fc39", x"5dc3e62e", x"f9bd0000", x"feab0000", x"cf080900", x"05560000", x"2c97007b", x"361db598", x"16d6024f", x"ed083c51"),
	(x"fb120000", x"49830000", x"75140a00", x"53ce0000", x"961a45a8", x"b65573ff", x"bf8a16d5", x"19fed62a", x"35a90000", x"5bc80000", x"95b10e80", x"3e060000", x"67471384", x"b1868180", x"7f954a8e", x"2752bbaf"),
	(x"37060000", x"ece00000", x"2fad0d80", x"689e0000", x"ddca5657", x"31ce47e7", x"d6c95e14", x"d3a451d4", x"b4370000", x"b79f0000", x"f3830c00", x"abf50000", x"3aee3b86", x"f972bd3c", x"99cfe8a3", x"a9350c55"),
	(x"ac480000", x"1ba60000", x"45fb1380", x"03430000", x"5a85316a", x"1fb250b6", x"fe72c7fe", x"91e478f6", x"1e4e0000", x"decf0000", x"6df80180", x"77240000", x"ec47079e", x"f4a0694e", x"cda31812", x"98aa496e"),
	(x"605c0000", x"bec50000", x"1f421400", x"38130000", x"11552295", x"982964ae", x"97318f3f", x"5bbeff08", x"9fd00000", x"32980000", x"0bca0300", x"e2d70000", x"b1ee2f9c", x"bc5455f2", x"2bf9ba3f", x"16cdfe94"),
	(x"2dd60000", x"f7f10000", x"23c91100", x"96b00000", x"072c1968", x"57466c0a", x"182865d3", x"1f83cf0c", x"53c40000", x"97fb0000", x"51730480", x"d9870000", x"fa3e3c63", x"3bcf61ea", x"42baf2fe", x"dc97796a"),
	(x"e1c20000", x"52920000", x"79701680", x"ade00000", x"4cfc0a97", x"d0dd5812", x"716b2d12", x"d5d948f2", x"d25a0000", x"7bac0000", x"37410600", x"4c740000", x"a7971461", x"733b5d56", x"a4e050d3", x"52f0ce90"),
	(x"d46b0000", x"095a0000", x"ecc11800", x"93e60000", x"2bbb1913", x"615bd992", x"0efe679c", x"f28bf35d", x"1ce10000", x"69e70000", x"d7e40280", x"21bc0000", x"56ca424d", x"74e8af29", x"64ff0c88", x"6c5ca315"),
	(x"187f0000", x"ac390000", x"b6781f80", x"a8b60000", x"606b0aec", x"e6c0ed8a", x"67bd2f5d", x"38d174a3", x"9d7f0000", x"85b00000", x"b1d60000", x"b44f0000", x"0b636a4f", x"3c1c9395", x"82a5aea5", x"e23b14ef"),
	(x"55f50000", x"e50d0000", x"8af31a80", x"06150000", x"76123111", x"29afe52e", x"e8a4c5b1", x"7cec44a7", x"516b0000", x"20d30000", x"eb6f0780", x"8f1f0000", x"40b379b0", x"bb87a78d", x"ebe6e664", x"28619311"),
	(x"99e10000", x"406e0000", x"d04a1d00", x"3d450000", x"3dc222ee", x"ae34d136", x"81e78d70", x"b6b6c359", x"d0f50000", x"cc840000", x"8d5d0500", x"1aec0000", x"1d1a51b2", x"f3739b31", x"0dbc4449", x"a60624eb"),
	(x"aee70000", x"ac8e0000", x"ffe71080", x"55db0000", x"e00874b9", x"9ffa96d1", x"572ed364", x"6512928d", x"64c20000", x"7b1b0000", x"7ede0900", x"b1190000", x"27f46a34", x"0a01260d", x"9473acea", x"0f3328be"),
	(x"62f30000", x"09ed0000", x"a55e1700", x"6e8b0000", x"abd86746", x"1861a2c9", x"3e6d9ba5", x"af481573", x"e55c0000", x"974c0000", x"18ec0b80", x"24ea0000", x"7a5d4236", x"42f51ab1", x"72290ec7", x"81549f44"),
	(x"2f790000", x"40d90000", x"99d51200", x"c0280000", x"bda15cbb", x"d70eaa6d", x"b1747149", x"eb752577", x"29480000", x"322f0000", x"42550c00", x"1fba0000", x"318d51c9", x"c56e2ea9", x"1b6a4606", x"4b0e18ba"),
	(x"e36d0000", x"e5ba0000", x"c36c1580", x"fb780000", x"f6714f44", x"50959e75", x"d8373988", x"212fa289", x"a8d60000", x"de780000", x"24670e80", x"8a490000", x"6c2479cb", x"8d9a1215", x"fd30e42b", x"c569af40"),
	(x"d6c40000", x"be720000", x"56dd1b00", x"c57e0000", x"91365cc0", x"e1131ff5", x"a7a27306", x"067d1926", x"666d0000", x"cc330000", x"c4c20a00", x"e7810000", x"9d792fe7", x"8a49e06a", x"3d2fb870", x"fbc5c2c5"),
	(x"1ad00000", x"1b110000", x"0c641c80", x"fe2e0000", x"dae64f3f", x"66882bed", x"cee13bc7", x"cc279ed8", x"e7f30000", x"20640000", x"a2f00880", x"72720000", x"c0d007e5", x"c2bddcd6", x"db751a5d", x"75a2753f"),
	(x"575a0000", x"52250000", x"30ef1980", x"508d0000", x"cc9f74c2", x"a9e72349", x"41f8d12b", x"881aaedc", x"2be70000", x"85070000", x"f8490f00", x"49220000", x"8b00141a", x"4526e8ce", x"b236529c", x"bff8f2c1"),
	(x"9b4e0000", x"f7460000", x"6a561e00", x"6bdd0000", x"874f673d", x"2e7c1751", x"28bb99ea", x"42402922", x"aa790000", x"69500000", x"9e7b0d80", x"dcd10000", x"d6a93c18", x"0dd2d472", x"546cf0b1", x"319f453b"),
	(x"1e4e0000", x"decf0000", x"6df80180", x"77240000", x"ec47079e", x"f4a0694e", x"cda31812", x"98aa496e", x"b2060000", x"c5690000", x"28031200", x"74670000", x"b6c236f4", x"eb1239f8", x"33d1dfec", x"094e3198"),
	(x"d25a0000", x"7bac0000", x"37410600", x"4c740000", x"a7971461", x"733b5d56", x"a4e050d3", x"52f0ce90", x"33980000", x"293e0000", x"4e311080", x"e1940000", x"eb6b1ef6", x"a3e60544", x"d58b7dc1", x"87298662"),
	(x"9fd00000", x"32980000", x"0bca0300", x"e2d70000", x"b1ee2f9c", x"bc5455f2", x"2bf9ba3f", x"16cdfe94", x"ff8c0000", x"8c5d0000", x"14881700", x"dac40000", x"a0bb0d09", x"247d315c", x"bcc83500", x"4d73019c"),
	(x"53c40000", x"97fb0000", x"51730480", x"d9870000", x"fa3e3c63", x"3bcf61ea", x"42baf2fe", x"dc97796a", x"7e120000", x"600a0000", x"72ba1580", x"4f370000", x"fd12250b", x"6c890de0", x"5a92972d", x"c314b666"),
	(x"666d0000", x"cc330000", x"c4c20a00", x"e7810000", x"9d792fe7", x"8a49e06a", x"3d2fb870", x"fbc5c2c5", x"b0a90000", x"72410000", x"921f1100", x"22ff0000", x"0c4f7327", x"6b5aff9f", x"9a8dcb76", x"fdb8dbe3"),
	(x"aa790000", x"69500000", x"9e7b0d80", x"dcd10000", x"d6a93c18", x"0dd2d472", x"546cf0b1", x"319f453b", x"31370000", x"9e160000", x"f42d1380", x"b70c0000", x"51e65b25", x"23aec323", x"7cd7695b", x"73df6c19"),
	(x"e7f30000", x"20640000", x"a2f00880", x"72720000", x"c0d007e5", x"c2bddcd6", x"db751a5d", x"75a2753f", x"fd230000", x"3b750000", x"ae941400", x"8c5c0000", x"1a3648da", x"a435f73b", x"1594219a", x"b985ebe7"),
	(x"2be70000", x"85070000", x"f8490f00", x"49220000", x"8b00141a", x"4526e8ce", x"b236529c", x"bff8f2c1", x"7cbd0000", x"d7220000", x"c8a61680", x"19af0000", x"479f60d8", x"ecc1cb87", x"f3ce83b7", x"37e25c1d"),
	(x"1ce10000", x"69e70000", x"d7e40280", x"21bc0000", x"56ca424d", x"74e8af29", x"64ff0c88", x"6c5ca315", x"c88a0000", x"60bd0000", x"3b251a80", x"b25a0000", x"7d715b5e", x"15b376bb", x"6a016b14", x"9ed75048"),
	(x"d0f50000", x"cc840000", x"8d5d0500", x"1aec0000", x"1d1a51b2", x"f3739b31", x"0dbc4449", x"a60624eb", x"49140000", x"8cea0000", x"5d171800", x"27a90000", x"20d8735c", x"5d474a07", x"8c5bc939", x"10b0e7b2"),
	(x"9d7f0000", x"85b00000", x"b1d60000", x"b44f0000", x"0b636a4f", x"3c1c9395", x"82a5aea5", x"e23b14ef", x"85000000", x"29890000", x"07ae1f80", x"1cf90000", x"6b0860a3", x"dadc7e1f", x"e51881f8", x"daea604c"),
	(x"516b0000", x"20d30000", x"eb6f0780", x"8f1f0000", x"40b379b0", x"bb87a78d", x"ebe6e664", x"28619311", x"049e0000", x"c5de0000", x"619c1d00", x"890a0000", x"36a148a1", x"922842a3", x"034223d5", x"548dd7b6"),
	(x"64c20000", x"7b1b0000", x"7ede0900", x"b1190000", x"27f46a34", x"0a01260d", x"9473acea", x"0f3328be", x"ca250000", x"d7950000", x"81391980", x"e4c20000", x"c7fc1e8d", x"95fbb0dc", x"c35d7f8e", x"6a21ba33"),
	(x"a8d60000", x"de780000", x"24670e80", x"8a490000", x"6c2479cb", x"8d9a1215", x"fd30e42b", x"c569af40", x"4bbb0000", x"3bc20000", x"e70b1b00", x"71310000", x"9a55368f", x"dd0f8c60", x"2507dda3", x"e4460dc9"),
	(x"e55c0000", x"974c0000", x"18ec0b80", x"24ea0000", x"7a5d4236", x"42f51ab1", x"72290ec7", x"81549f44", x"87af0000", x"9ea10000", x"bdb21c80", x"4a610000", x"d1852570", x"5a94b878", x"4c449562", x"2e1c8a37"),
	(x"29480000", x"322f0000", x"42550c00", x"1fba0000", x"318d51c9", x"c56e2ea9", x"1b6a4606", x"4b0e18ba", x"06310000", x"72f60000", x"db801e00", x"df920000", x"8c2c0d72", x"126084c4", x"aa1e374f", x"a07b3dcd"),
	(x"b2060000", x"c5690000", x"28031200", x"74670000", x"b6c236f4", x"eb1239f8", x"33d1dfec", x"094e3198", x"ac480000", x"1ba60000", x"45fb1380", x"03430000", x"5a85316a", x"1fb250b6", x"fe72c7fe", x"91e478f6"),
	(x"7e120000", x"600a0000", x"72ba1580", x"4f370000", x"fd12250b", x"6c890de0", x"5a92972d", x"c314b666", x"2dd60000", x"f7f10000", x"23c91100", x"96b00000", x"072c1968", x"57466c0a", x"182865d3", x"1f83cf0c"),
	(x"33980000", x"293e0000", x"4e311080", x"e1940000", x"eb6b1ef6", x"a3e60544", x"d58b7dc1", x"87298662", x"e1c20000", x"52920000", x"79701680", x"ade00000", x"4cfc0a97", x"d0dd5812", x"716b2d12", x"d5d948f2"),
	(x"ff8c0000", x"8c5d0000", x"14881700", x"dac40000", x"a0bb0d09", x"247d315c", x"bcc83500", x"4d73019c", x"605c0000", x"bec50000", x"1f421400", x"38130000", x"11552295", x"982964ae", x"97318f3f", x"5bbeff08"),
	(x"ca250000", x"d7950000", x"81391980", x"e4c20000", x"c7fc1e8d", x"95fbb0dc", x"c35d7f8e", x"6a21ba33", x"aee70000", x"ac8e0000", x"ffe71080", x"55db0000", x"e00874b9", x"9ffa96d1", x"572ed364", x"6512928d"),
	(x"06310000", x"72f60000", x"db801e00", x"df920000", x"8c2c0d72", x"126084c4", x"aa1e374f", x"a07b3dcd", x"2f790000", x"40d90000", x"99d51200", x"c0280000", x"bda15cbb", x"d70eaa6d", x"b1747149", x"eb752577"),
	(x"4bbb0000", x"3bc20000", x"e70b1b00", x"71310000", x"9a55368f", x"dd0f8c60", x"2507dda3", x"e4460dc9", x"e36d0000", x"e5ba0000", x"c36c1580", x"fb780000", x"f6714f44", x"50959e75", x"d8373988", x"212fa289"),
	(x"87af0000", x"9ea10000", x"bdb21c80", x"4a610000", x"d1852570", x"5a94b878", x"4c449562", x"2e1c8a37", x"62f30000", x"09ed0000", x"a55e1700", x"6e8b0000", x"abd86746", x"1861a2c9", x"3e6d9ba5", x"af481573"),
	(x"b0a90000", x"72410000", x"921f1100", x"22ff0000", x"0c4f7327", x"6b5aff9f", x"9a8dcb76", x"fdb8dbe3", x"d6c40000", x"be720000", x"56dd1b00", x"c57e0000", x"91365cc0", x"e1131ff5", x"a7a27306", x"067d1926"),
	(x"7cbd0000", x"d7220000", x"c8a61680", x"19af0000", x"479f60d8", x"ecc1cb87", x"f3ce83b7", x"37e25c1d", x"575a0000", x"52250000", x"30ef1980", x"508d0000", x"cc9f74c2", x"a9e72349", x"41f8d12b", x"881aaedc"),
	(x"31370000", x"9e160000", x"f42d1380", x"b70c0000", x"51e65b25", x"23aec323", x"7cd7695b", x"73df6c19", x"9b4e0000", x"f7460000", x"6a561e00", x"6bdd0000", x"874f673d", x"2e7c1751", x"28bb99ea", x"42402922"),
	(x"fd230000", x"3b750000", x"ae941400", x"8c5c0000", x"1a3648da", x"a435f73b", x"1594219a", x"b985ebe7", x"1ad00000", x"1b110000", x"0c641c80", x"fe2e0000", x"dae64f3f", x"66882bed", x"cee13bc7", x"cc279ed8"),
	(x"c88a0000", x"60bd0000", x"3b251a80", x"b25a0000", x"7d715b5e", x"15b376bb", x"6a016b14", x"9ed75048", x"d46b0000", x"095a0000", x"ecc11800", x"93e60000", x"2bbb1913", x"615bd992", x"0efe679c", x"f28bf35d"),
	(x"049e0000", x"c5de0000", x"619c1d00", x"890a0000", x"36a148a1", x"922842a3", x"034223d5", x"548dd7b6", x"55f50000", x"e50d0000", x"8af31a80", x"06150000", x"76123111", x"29afe52e", x"e8a4c5b1", x"7cec44a7"),
	(x"49140000", x"8cea0000", x"5d171800", x"27a90000", x"20d8735c", x"5d474a07", x"8c5bc939", x"10b0e7b2", x"99e10000", x"406e0000", x"d04a1d00", x"3d450000", x"3dc222ee", x"ae34d136", x"81e78d70", x"b6b6c359"),
	(x"85000000", x"29890000", x"07ae1f80", x"1cf90000", x"6b0860a3", x"dadc7e1f", x"e51881f8", x"daea604c", x"187f0000", x"ac390000", x"b6781f80", x"a8b60000", x"606b0aec", x"e6c0ed8a", x"67bd2f5d", x"38d174a3"),
	(x"aec30000", x"9c4f0001", x"79d1e000", x"2c150000", x"45cc75b3", x"6650b736", x"ab92f78f", x"a312567b", x"db250000", x"09290000", x"49aac000", x"81e10000", x"cafe6b59", x"42793431", x"43566b76", x"e86cba2e"),
	(x"62d70000", x"392c0001", x"2368e780", x"17450000", x"0e1c664c", x"e1cb832e", x"c2d1bf4e", x"6948d185", x"5abb0000", x"e57e0000", x"2f98c280", x"14120000", x"9757435b", x"0a8d088d", x"a50cc95b", x"660b0dd4"),
	(x"2f5d0000", x"70180001", x"1fe3e280", x"b9e60000", x"18655db1", x"2ea48b8a", x"4dc855a2", x"2d75e181", x"96af0000", x"401d0000", x"7521c500", x"2f420000", x"dc8750a4", x"8d163c95", x"cc4f819a", x"ac518a2a"),
	(x"e3490000", x"d57b0001", x"455ae500", x"82b60000", x"53b54e4e", x"a93fbf92", x"248b1d63", x"e72f667f", x"17310000", x"ac4a0000", x"1313c780", x"bab10000", x"812e78a6", x"c5e20029", x"2a1523b7", x"22363dd0"),
	(x"d6e00000", x"8eb30001", x"d0ebeb80", x"bcb00000", x"34f25dca", x"18b93e12", x"5b1e57ed", x"c07dddd0", x"d98a0000", x"be010000", x"f3b6c300", x"d7790000", x"70732e8a", x"c231f256", x"ea0a7fec", x"1c9a5055"),
	(x"1af40000", x"2bd00001", x"8a52ec00", x"87e00000", x"7f224e35", x"9f220a0a", x"325d1f2c", x"0a275a2e", x"58140000", x"52560000", x"9584c180", x"428a0000", x"2dda0688", x"8ac5ceea", x"0c50ddc1", x"92fde7af"),
	(x"577e0000", x"62e40001", x"b6d9e900", x"29430000", x"695b75c8", x"504d02ae", x"bd44f5c0", x"4e1a6a2a", x"94000000", x"f7350000", x"cf3dc600", x"79da0000", x"660a1577", x"0d5efaf2", x"65139500", x"58a76051"),
	(x"9b6a0000", x"c7870001", x"ec60ee80", x"12130000", x"228b6637", x"d7d636b6", x"d407bd01", x"8440edd4", x"159e0000", x"1b620000", x"a90fc480", x"ec290000", x"3ba33d75", x"45aac64e", x"8349372d", x"d6c0d7ab"),
	(x"ac6c0000", x"2b670001", x"c3cde300", x"7a8d0000", x"ff413060", x"e6187151", x"02cee315", x"57e4bc00", x"a1a90000", x"acfd0000", x"5a8cc880", x"47dc0000", x"014d06f3", x"bcd87b72", x"1a86df8e", x"7ff5dbfe"),
	(x"60780000", x"8e040001", x"9974e480", x"41dd0000", x"b491239f", x"61834549", x"6b8dabd4", x"9dbe3bfe", x"20370000", x"40aa0000", x"3cbeca00", x"d22f0000", x"5ce42ef1", x"f42c47ce", x"fcdc7da3", x"f1926c04"),
	(x"2df20000", x"c7300001", x"a5ffe180", x"ef7e0000", x"a2e81862", x"aeec4ded", x"e4944138", x"d9830bfa", x"ec230000", x"e5c90000", x"6607cd80", x"e97f0000", x"17343d0e", x"73b773d6", x"959f3562", x"3bc8ebfa"),
	(x"e1e60000", x"62530001", x"ff46e600", x"d42e0000", x"e9380b9d", x"297779f5", x"8dd709f9", x"13d98c04", x"6dbd0000", x"099e0000", x"0035cf00", x"7c8c0000", x"4a9d150c", x"3b434f6a", x"73c5974f", x"b5af5c00"),
	(x"d44f0000", x"399b0001", x"6af7e880", x"ea280000", x"8e7f1819", x"98f1f875", x"f2424377", x"348b37ab", x"a3060000", x"1bd50000", x"e090cb80", x"11440000", x"bbc04320", x"3c90bd15", x"b3dacb14", x"8b033185"),
	(x"185b0000", x"9cf80001", x"304eef00", x"d1780000", x"c5af0be6", x"1f6acc6d", x"9b010bb6", x"fed1b055", x"22980000", x"f7820000", x"86a2c900", x"84b70000", x"e6696b22", x"746481a9", x"55806939", x"0564867f"),
	(x"55d10000", x"d5cc0001", x"0cc5ea00", x"7fdb0000", x"d3d6301b", x"d005c4c9", x"1418e15a", x"baec8051", x"ee8c0000", x"52e10000", x"dc1bce80", x"bfe70000", x"adb978dd", x"f3ffb5b1", x"3cc321f8", x"cf3e0181"),
	(x"99c50000", x"70af0001", x"567ced80", x"448b0000", x"980623e4", x"579ef0d1", x"7d5ba99b", x"70b607af", x"6f120000", x"beb60000", x"ba29cc00", x"2a140000", x"f01050df", x"bb0b890d", x"da9983d5", x"4159b67b"),
	(x"028b0000", x"87e90001", x"3c2af380", x"2f560000", x"1f4944d9", x"79e2e780", x"55e03071", x"32f62e8d", x"c56b0000", x"d7e60000", x"2452c180", x"f6c50000", x"26b96cc7", x"b6d95d7f", x"8ef57364", x"70c6f340"),
	(x"ce9f0000", x"228a0001", x"6693f400", x"14060000", x"54995726", x"fe79d398", x"3ca378b0", x"f8aca973", x"44f50000", x"3bb10000", x"4260c300", x"63360000", x"7b1044c5", x"fe2d61c3", x"68afd149", x"fea144ba"),
	(x"83150000", x"6bbe0001", x"5a18f100", x"baa50000", x"42e06cdb", x"3116db3c", x"b3ba925c", x"bc919977", x"88e10000", x"9ed20000", x"18d9c480", x"58660000", x"30c0573a", x"79b655db", x"01ec9988", x"34fbc344"),
	(x"4f010000", x"cedd0001", x"00a1f680", x"81f50000", x"09307f24", x"b68def24", x"daf9da9d", x"76cb1e89", x"097f0000", x"72850000", x"7eebc600", x"cd950000", x"6d697f38", x"31426967", x"e7b63ba5", x"ba9c74be"),
	(x"7aa80000", x"95150001", x"9510f800", x"bff30000", x"6e776ca0", x"070b6ea4", x"a56c9013", x"5199a526", x"c7c40000", x"60ce0000", x"9e4ec280", x"a05d0000", x"9c342914", x"36919b18", x"27a967fe", x"8430193b"),
	(x"b6bc0000", x"30760001", x"cfa9ff80", x"84a30000", x"25a77f5f", x"80905abc", x"cc2fd8d2", x"9bc322d8", x"465a0000", x"8c990000", x"f87cc000", x"35ae0000", x"c19d0116", x"7e65a7a4", x"c1f3c5d3", x"0a57aec1"),
	(x"fb360000", x"79420001", x"f322fa80", x"2a000000", x"33de44a2", x"4fff5218", x"4336323e", x"dffe12dc", x"8a4e0000", x"29fa0000", x"a2c5c780", x"0efe0000", x"8a4d12e9", x"f9fe93bc", x"a8b08d12", x"c00d293f"),
	(x"37220000", x"dc210001", x"a99bfd00", x"11500000", x"780e575d", x"c8646600", x"2a757aff", x"15a49522", x"0bd00000", x"c5ad0000", x"c4f7c500", x"9b0d0000", x"d7e43aeb", x"b10aaf00", x"4eea2f3f", x"4e6a9ec5"),
	(x"00240000", x"30c10001", x"8636f080", x"79ce0000", x"a5c4010a", x"f9aa21e7", x"fcbc24eb", x"c600c4f6", x"bfe70000", x"72320000", x"3774c900", x"30f80000", x"ed0a016d", x"4878123c", x"d725c79c", x"e75f9290"),
	(x"cc300000", x"95a20001", x"dc8ff700", x"429e0000", x"ee1412f5", x"7e3115ff", x"95ff6c2a", x"0c5a4308", x"3e790000", x"9e650000", x"5146cb80", x"a50b0000", x"b0a3296f", x"008c2e80", x"317f65b1", x"6938256a"),
	(x"81ba0000", x"dc960001", x"e004f200", x"ec3d0000", x"f86d2908", x"b15e1d5b", x"1ae686c6", x"4867730c", x"f26d0000", x"3b060000", x"0bffcc00", x"9e5b0000", x"fb733a90", x"87171a98", x"583c2d70", x"a362a294"),
	(x"4dae0000", x"79f50001", x"babdf580", x"d76d0000", x"b3bd3af7", x"36c52943", x"73a5ce07", x"823df4f2", x"73f30000", x"d7510000", x"6dcdce80", x"0ba80000", x"a6da1292", x"cfe32624", x"be668f5d", x"2d05156e"),
	(x"78070000", x"223d0001", x"2f0cfb00", x"e96b0000", x"d4fa2973", x"8743a8c3", x"0c308489", x"a56f4f5d", x"bd480000", x"c51a0000", x"8d68ca00", x"66600000", x"578744be", x"c830d45b", x"7e79d306", x"13a978eb"),
	(x"b4130000", x"875e0001", x"75b5fc80", x"d23b0000", x"9f2a3a8c", x"00d89cdb", x"6573cc48", x"6f35c8a3", x"3cd60000", x"294d0000", x"eb5ac880", x"f3930000", x"0a2e6cbc", x"80c4e8e7", x"9823712b", x"9dcecf11"),
	(x"f9990000", x"ce6a0001", x"493ef980", x"7c980000", x"89530171", x"cfb7947f", x"ea6a26a4", x"2b08f8a7", x"f0c20000", x"8c2e0000", x"b1e3cf00", x"c8c30000", x"41fe7f43", x"075fdcff", x"f16039ea", x"579448ef"),
	(x"358d0000", x"6b090001", x"1387fe00", x"47c80000", x"c283128e", x"482ca067", x"83296e65", x"e1527f59", x"715c0000", x"60790000", x"d7d1cd80", x"5d300000", x"1c575741", x"4fabe043", x"173a9bc7", x"d9f3ff15"),
	(x"b08d0000", x"42800001", x"1429e180", x"5b310000", x"a98b722d", x"92f0de78", x"6631ef9d", x"3bb81f15", x"69230000", x"cc400000", x"61a9d200", x"f5860000", x"7c3c5dad", x"a96b0dc9", x"7087b49a", x"e1228bb6"),
	(x"7c990000", x"e7e30001", x"4e90e600", x"60610000", x"e25b61d2", x"156bea60", x"0f72a75c", x"f1e298eb", x"e8bd0000", x"20170000", x"079bd080", x"60750000", x"219575af", x"e19f3175", x"96dd16b7", x"6f453c4c"),
	(x"31130000", x"aed70001", x"721be300", x"cec20000", x"f4225a2f", x"da04e2c4", x"806b4db0", x"b5dfa8ef", x"24a90000", x"85740000", x"5d22d700", x"5b250000", x"6a456650", x"6604056d", x"ff9e5e76", x"a51fbbb2"),
	(x"fd070000", x"0bb40001", x"28a2e480", x"f5920000", x"bff249d0", x"5d9fd6dc", x"e9280571", x"7f852f11", x"a5370000", x"69230000", x"3b10d580", x"ced60000", x"37ec4e52", x"2ef039d1", x"19c4fc5b", x"2b780c48"),
	(x"c8ae0000", x"507c0001", x"bd13ea00", x"cb940000", x"d8b55a54", x"ec19575c", x"96bd4fff", x"58d794be", x"6b8c0000", x"7b680000", x"dbb5d100", x"a31e0000", x"c6b1187e", x"2923cbae", x"d9dba000", x"15d461cd"),
	(x"04ba0000", x"f51f0001", x"e7aaed80", x"f0c40000", x"936549ab", x"6b826344", x"fffe073e", x"928d1340", x"ea120000", x"973f0000", x"bd87d380", x"36ed0000", x"9b18307c", x"61d7f712", x"3f81022d", x"9bb3d637"),
	(x"49300000", x"bc2b0001", x"db21e880", x"5e670000", x"851c7256", x"a4ed6be0", x"70e7edd2", x"d6b02344", x"26060000", x"325c0000", x"e73ed400", x"0dbd0000", x"d0c82383", x"e64cc30a", x"56c24aec", x"51e951c9"),
	(x"85240000", x"19480001", x"8198ef00", x"65370000", x"cecc61a9", x"23765ff8", x"19a4a513", x"1ceaa4ba", x"a7980000", x"de0b0000", x"810cd680", x"984e0000", x"8d610b81", x"aeb8ffb6", x"b098e8c1", x"df8ee633"),
	(x"b2220000", x"f5a80001", x"ae35e280", x"0da90000", x"130637fe", x"12b8181f", x"cf6dfb07", x"cf4ef56e", x"13af0000", x"69940000", x"728fda80", x"33bb0000", x"b78f3007", x"57ca428a", x"29570062", x"76bbea66"),
	(x"7e360000", x"50cb0001", x"f48ce500", x"36f90000", x"58d62401", x"95232c07", x"a62eb3c6", x"05147290", x"92310000", x"85c30000", x"14bdd800", x"a6480000", x"ea261805", x"1f3e7e36", x"cf0da24f", x"f8dc5d9c"),
	(x"33bc0000", x"19ff0001", x"c807e000", x"985a0000", x"4eaf1ffc", x"5a4c24a3", x"2937592a", x"41294294", x"5e250000", x"20a00000", x"4e04df80", x"9d180000", x"a1f60bfa", x"98a54a2e", x"a64eea8e", x"3286da62"),
	(x"ffa80000", x"bc9c0001", x"92bee780", x"a30a0000", x"057f0c03", x"ddd710bb", x"407411eb", x"8b73c56a", x"dfbb0000", x"ccf70000", x"2836dd00", x"08eb0000", x"fc5f23f8", x"d0517692", x"401448a3", x"bce16d98"),
	(x"ca010000", x"e7540001", x"070fe900", x"9d0c0000", x"62381f87", x"6c51913b", x"3fe15b65", x"ac217ec5", x"11000000", x"debc0000", x"c893d980", x"65230000", x"0d0275d4", x"d78284ed", x"800b14f8", x"824d001d"),
	(x"06150000", x"42370001", x"5db6ee80", x"a65c0000", x"29e80c78", x"ebcaa523", x"56a213a4", x"667bf93b", x"909e0000", x"32eb0000", x"aea1db00", x"f0d00000", x"50ab5dd6", x"9f76b851", x"6651b6d5", x"0c2ab7e7"),
	(x"4b9f0000", x"0b030001", x"613deb80", x"08ff0000", x"3f913785", x"24a5ad87", x"d9bbf948", x"2246c93f", x"5c8a0000", x"97880000", x"f418dc80", x"cb800000", x"1b7b4e29", x"18ed8c49", x"0f12fe14", x"c6703019"),
	(x"878b0000", x"ae600001", x"3b84ec00", x"33af0000", x"7441247a", x"a33e999f", x"b0f8b189", x"e81c4ec1", x"dd140000", x"7bdf0000", x"922ade00", x"5e730000", x"46d2662b", x"5019b0f5", x"e9485c39", x"481787e3"),
	(x"1cc50000", x"59260001", x"51d2f200", x"58720000", x"f30e4347", x"8d428ece", x"98432863", x"aa5c67e3", x"776d0000", x"128f0000", x"0c51d380", x"82a20000", x"907b5a33", x"5dcb6487", x"bd24ac88", x"7988c2d8"),
	(x"d0d10000", x"fc450001", x"0b6bf580", x"63220000", x"b8de50b8", x"0ad9bad6", x"f10060a2", x"6006e01d", x"f6f30000", x"fed80000", x"6a63d100", x"17510000", x"cdd27231", x"153f583b", x"5b7e0ea5", x"f7ef7522"),
	(x"9d5b0000", x"b5710001", x"37e0f080", x"cd810000", x"aea76b45", x"c5b6b272", x"7e198a4e", x"243bd019", x"3ae70000", x"5bbb0000", x"30dad680", x"2c010000", x"860261ce", x"92a46c23", x"323d4664", x"3db5f2dc"),
	(x"514f0000", x"10120001", x"6d59f700", x"f6d10000", x"e57778ba", x"422d866a", x"175ac28f", x"ee6157e7", x"bb790000", x"b7ec0000", x"56e8d400", x"b9f20000", x"dbab49cc", x"da50509f", x"d467e449", x"b3d24526"),
	(x"64e60000", x"4bda0001", x"f8e8f980", x"c8d70000", x"82306b3e", x"f3ab07ea", x"68cf8801", x"c933ec48", x"75c20000", x"a5a70000", x"b64dd080", x"d43a0000", x"2af61fe0", x"dd83a2e0", x"1478b812", x"8d7e28a3"),
	(x"a8f20000", x"eeb90001", x"a251fe00", x"f3870000", x"c9e078c1", x"743033f2", x"018cc0c0", x"03696bb6", x"f45c0000", x"49f00000", x"d07fd200", x"41c90000", x"775f37e2", x"95779e5c", x"f2221a3f", x"03199f59"),
	(x"e5780000", x"a78d0001", x"9edafb00", x"5d240000", x"df99433c", x"bb5f3b56", x"8e952a2c", x"47545bb2", x"38480000", x"ec930000", x"8ac6d580", x"7a990000", x"3c8f241d", x"12ecaa44", x"9b6152fe", x"c94318a7"),
	(x"296c0000", x"02ee0001", x"c463fc80", x"66740000", x"944950c3", x"3cc40f4e", x"e7d662ed", x"8d0edc4c", x"b9d60000", x"00c40000", x"ecf4d700", x"ef6a0000", x"61260c1f", x"5a1896f8", x"7d3bf0d3", x"4724af5d"),
	(x"1e6a0000", x"ee0e0001", x"ebcef100", x"0eea0000", x"49830694", x"0d0a48a9", x"311f3cf9", x"5eaa8d98", x"0de10000", x"b75b0000", x"1f77db00", x"449f0000", x"5bc83799", x"a36a2bc4", x"e4f41870", x"ee11a308"),
	(x"d27e0000", x"4b6d0001", x"b177f680", x"35ba0000", x"0253156b", x"8a917cb1", x"585c7438", x"94f00a66", x"8c7f0000", x"5b0c0000", x"7945d980", x"d16c0000", x"06611f9b", x"eb9e1778", x"02aeba5d", x"607614f2"),
	(x"9ff40000", x"02590001", x"8dfcf380", x"9b190000", x"142a2e96", x"45fe7415", x"d7459ed4", x"d0cd3a62", x"406b0000", x"fe6f0000", x"23fcde00", x"ea3c0000", x"4db10c64", x"6c052360", x"6bedf29c", x"aa2c930c"),
	(x"53e00000", x"a73a0001", x"d745f400", x"a0490000", x"5ffa3d69", x"c265400d", x"be06d615", x"1a97bd9c", x"c1f50000", x"12380000", x"45cedc80", x"7fcf0000", x"10182466", x"24f11fdc", x"8db750b1", x"244b24f6"),
	(x"66490000", x"fcf20001", x"42f4fa80", x"9e4f0000", x"38bd2eed", x"73e3c18d", x"c1939c9b", x"3dc50633", x"0f4e0000", x"00730000", x"a56bd800", x"12070000", x"e145724a", x"2322eda3", x"4da80cea", x"1ae74973"),
	(x"aa5d0000", x"59910001", x"184dfd00", x"a51f0000", x"736d3d12", x"f478f595", x"a8d0d45a", x"f79f81cd", x"8ed00000", x"ec240000", x"c359da80", x"87f40000", x"bcec5a48", x"6bd6d11f", x"abf2aec7", x"9480fe89"),
	(x"e7d70000", x"10a50001", x"24c6f800", x"0bbc0000", x"651406ef", x"3b17fd31", x"27c93eb6", x"b3a2b1c9", x"42c40000", x"49470000", x"99e0dd00", x"bca40000", x"f73c49b7", x"ec4de507", x"c2b1e606", x"5eda7977"),
	(x"2bc30000", x"b5c60001", x"7e7fff80", x"30ec0000", x"2ec41510", x"bc8cc929", x"4e8a7677", x"79f83637", x"c35a0000", x"a5100000", x"ffd2df80", x"29570000", x"aa9561b5", x"a4b9d9bb", x"24eb442b", x"d0bdce8d"),
	(x"db250000", x"09290000", x"49aac000", x"81e10000", x"cafe6b59", x"42793431", x"43566b76", x"e86cba2e", x"75e60000", x"95660001", x"307b2000", x"adf40000", x"8f321eea", x"24298307", x"e8c49cf9", x"4b7eec55"),
	(x"17310000", x"ac4a0000", x"1313c780", x"bab10000", x"812e78a6", x"c5e20029", x"2a1523b7", x"22363dd0", x"f4780000", x"79310001", x"56492280", x"38070000", x"d29b36e8", x"6cddbfbb", x"0e9e3ed4", x"c5195baf"),
	(x"5abb0000", x"e57e0000", x"2f98c280", x"14120000", x"9757435b", x"0a8d088d", x"a50cc95b", x"660b0dd4", x"386c0000", x"dc520001", x"0cf02500", x"03570000", x"994b2517", x"eb468ba3", x"67dd7615", x"0f43dc51"),
	(x"96af0000", x"401d0000", x"7521c500", x"2f420000", x"dc8750a4", x"8d163c95", x"cc4f819a", x"ac518a2a", x"b9f20000", x"30050001", x"6ac22780", x"96a40000", x"c4e20d15", x"a3b2b71f", x"8187d438", x"81246bab"),
	(x"a3060000", x"1bd50000", x"e090cb80", x"11440000", x"bbc04320", x"3c90bd15", x"b3dacb14", x"8b033185", x"77490000", x"224e0001", x"8a672300", x"fb6c0000", x"35bf5b39", x"a4614560", x"41988863", x"bf88062e"),
	(x"6f120000", x"beb60000", x"ba29cc00", x"2a140000", x"f01050df", x"bb0b890d", x"da9983d5", x"4159b67b", x"f6d70000", x"ce190001", x"ec552180", x"6e9f0000", x"6816733b", x"ec9579dc", x"a7c22a4e", x"31efb1d4"),
	(x"22980000", x"f7820000", x"86a2c900", x"84b70000", x"e6696b22", x"746481a9", x"55806939", x"0564867f", x"3ac30000", x"6b7a0001", x"b6ec2600", x"55cf0000", x"23c660c4", x"6b0e4dc4", x"ce81628f", x"fbb5362a"),
	(x"ee8c0000", x"52e10000", x"dc1bce80", x"bfe70000", x"adb978dd", x"f3ffb5b1", x"3cc321f8", x"cf3e0181", x"bb5d0000", x"872d0001", x"d0de2480", x"c03c0000", x"7e6f48c6", x"23fa7178", x"28dbc0a2", x"75d281d0"),
	(x"d98a0000", x"be010000", x"f3b6c300", x"d7790000", x"70732e8a", x"c231f256", x"ea0a7fec", x"1c9a5055", x"0f6a0000", x"30b20001", x"235d2880", x"6bc90000", x"44817340", x"da88cc44", x"b1142801", x"dce78d85"),
	(x"159e0000", x"1b620000", x"a90fc480", x"ec290000", x"3ba33d75", x"45aac64e", x"8349372d", x"d6c0d7ab", x"8ef40000", x"dce50001", x"456f2a00", x"fe3a0000", x"19285b42", x"927cf0f8", x"574e8a2c", x"52803a7f"),
	(x"58140000", x"52560000", x"9584c180", x"428a0000", x"2dda0688", x"8ac5ceea", x"0c50ddc1", x"92fde7af", x"42e00000", x"79860001", x"1fd62d80", x"c56a0000", x"52f848bd", x"15e7c4e0", x"3e0dc2ed", x"98dabd81"),
	(x"94000000", x"f7350000", x"cf3dc600", x"79da0000", x"660a1577", x"0d5efaf2", x"65139500", x"58a76051", x"c37e0000", x"95d10001", x"79e42f00", x"50990000", x"0f5160bf", x"5d13f85c", x"d85760c0", x"16bd0a7b"),
	(x"a1a90000", x"acfd0000", x"5a8cc880", x"47dc0000", x"014d06f3", x"bcd87b72", x"1a86df8e", x"7ff5dbfe", x"0dc50000", x"879a0001", x"99412b80", x"3d510000", x"fe0c3693", x"5ac00a23", x"18483c9b", x"281167fe"),
	(x"6dbd0000", x"099e0000", x"0035cf00", x"7c8c0000", x"4a9d150c", x"3b434f6a", x"73c5974f", x"b5af5c00", x"8c5b0000", x"6bcd0001", x"ff732900", x"a8a20000", x"a3a51e91", x"1234369f", x"fe129eb6", x"a676d004"),
	(x"20370000", x"40aa0000", x"3cbeca00", x"d22f0000", x"5ce42ef1", x"f42c47ce", x"fcdc7da3", x"f1926c04", x"404f0000", x"ceae0001", x"a5ca2e80", x"93f20000", x"e8750d6e", x"95af0287", x"9751d677", x"6c2c57fa"),
	(x"ec230000", x"e5c90000", x"6607cd80", x"e97f0000", x"17343d0e", x"73b773d6", x"959f3562", x"3bc8ebfa", x"c1d10000", x"22f90001", x"c3f82c00", x"06010000", x"b5dc256c", x"dd5b3e3b", x"710b745a", x"e24be000"),
	(x"776d0000", x"128f0000", x"0c51d380", x"82a20000", x"907b5a33", x"5dcb6487", x"bd24ac88", x"7988c2d8", x"6ba80000", x"4ba90001", x"5d832180", x"dad00000", x"63751974", x"d089ea49", x"256784eb", x"d3d4a53b"),
	(x"bb790000", x"b7ec0000", x"56e8d400", x"b9f20000", x"dbab49cc", x"da50509f", x"d467e449", x"b3d24526", x"ea360000", x"a7fe0001", x"3bb12300", x"4f230000", x"3edc3176", x"987dd6f5", x"c33d26c6", x"5db312c1"),
	(x"f6f30000", x"fed80000", x"6a63d100", x"17510000", x"cdd27231", x"153f583b", x"5b7e0ea5", x"f7ef7522", x"26220000", x"029d0001", x"61082480", x"74730000", x"750c2289", x"1fe6e2ed", x"aa7e6e07", x"97e9953f"),
	(x"3ae70000", x"5bbb0000", x"30dad680", x"2c010000", x"860261ce", x"92a46c23", x"323d4664", x"3db5f2dc", x"a7bc0000", x"eeca0001", x"073a2600", x"e1800000", x"28a50a8b", x"5712de51", x"4c24cc2a", x"198e22c5"),
	(x"0f4e0000", x"00730000", x"a56bd800", x"12070000", x"e145724a", x"2322eda3", x"4da80cea", x"1ae74973", x"69070000", x"fc810001", x"e79f2280", x"8c480000", x"d9f85ca7", x"50c12c2e", x"8c3b9071", x"27224f40"),
	(x"c35a0000", x"a5100000", x"ffd2df80", x"29570000", x"aa9561b5", x"a4b9d9bb", x"24eb442b", x"d0bdce8d", x"e8990000", x"10d60001", x"81ad2000", x"19bb0000", x"845174a5", x"18351092", x"6a61325c", x"a945f8ba"),
	(x"8ed00000", x"ec240000", x"c359da80", x"87f40000", x"bcec5a48", x"6bd6d11f", x"abf2aec7", x"9480fe89", x"248d0000", x"b5b50001", x"db142780", x"22eb0000", x"cf81675a", x"9fae248a", x"03227a9d", x"631f7f44"),
	(x"42c40000", x"49470000", x"99e0dd00", x"bca40000", x"f73c49b7", x"ec4de507", x"c2b1e606", x"5eda7977", x"a5130000", x"59e20001", x"bd262500", x"b7180000", x"92284f58", x"d75a1836", x"e578d8b0", x"ed78c8be"),
	(x"75c20000", x"a5a70000", x"b64dd080", x"d43a0000", x"2af61fe0", x"dd83a2e0", x"1478b812", x"8d7e28a3", x"11240000", x"ee7d0001", x"4ea52900", x"1ced0000", x"a8c674de", x"2e28a50a", x"7cb73013", x"444dc4eb"),
	(x"b9d60000", x"00c40000", x"ecf4d700", x"ef6a0000", x"61260c1f", x"5a1896f8", x"7d3bf0d3", x"4724af5d", x"90ba0000", x"022a0001", x"28972b80", x"891e0000", x"f56f5cdc", x"66dc99b6", x"9aed923e", x"ca2a7311"),
	(x"f45c0000", x"49f00000", x"d07fd200", x"41c90000", x"775f37e2", x"95779e5c", x"f2221a3f", x"03199f59", x"5cae0000", x"a7490001", x"722e2c00", x"b24e0000", x"bebf4f23", x"e147adae", x"f3aedaff", x"0070f4ef"),
	(x"38480000", x"ec930000", x"8ac6d580", x"7a990000", x"3c8f241d", x"12ecaa44", x"9b6152fe", x"c94318a7", x"dd300000", x"4b1e0001", x"141c2e80", x"27bd0000", x"e3166721", x"a9b39112", x"15f478d2", x"8e174315"),
	(x"0de10000", x"b75b0000", x"1f77db00", x"449f0000", x"5bc83799", x"a36a2bc4", x"e4f41870", x"ee11a308", x"138b0000", x"59550001", x"f4b92a00", x"4a750000", x"124b310d", x"ae60636d", x"d5eb2489", x"b0bb2e90"),
	(x"c1f50000", x"12380000", x"45cedc80", x"7fcf0000", x"10182466", x"24f11fdc", x"8db750b1", x"244b24f6", x"92150000", x"b5020001", x"928b2880", x"df860000", x"4fe2190f", x"e6945fd1", x"33b186a4", x"3edc996a"),
	(x"8c7f0000", x"5b0c0000", x"7945d980", x"d16c0000", x"06611f9b", x"eb9e1778", x"02aeba5d", x"607614f2", x"5e010000", x"10610001", x"c8322f00", x"e4d60000", x"04320af0", x"610f6bc9", x"5af2ce65", x"f4861e94"),
	(x"406b0000", x"fe6f0000", x"23fcde00", x"ea3c0000", x"4db10c64", x"6c052360", x"6bedf29c", x"aa2c930c", x"df9f0000", x"fc360001", x"ae002d80", x"71250000", x"599b22f2", x"29fb5775", x"bca86c48", x"7ae1a96e"),
	(x"c56b0000", x"d7e60000", x"2452c180", x"f6c50000", x"26b96cc7", x"b6d95d7f", x"8ef57364", x"70c6f340", x"c7e00000", x"500f0001", x"18783200", x"d9930000", x"39f0281e", x"cf3bbaff", x"db154315", x"4230ddcd"),
	(x"097f0000", x"72850000", x"7eebc600", x"cd950000", x"6d697f38", x"31426967", x"e7b63ba5", x"ba9c74be", x"467e0000", x"bc580001", x"7e4a3080", x"4c600000", x"6459001c", x"87cf8643", x"3d4fe138", x"cc576a37"),
	(x"44f50000", x"3bb10000", x"4260c300", x"63360000", x"7b1044c5", x"fe2d61c3", x"68afd149", x"fea144ba", x"8a6a0000", x"193b0001", x"24f33700", x"77300000", x"2f8913e3", x"0054b25b", x"540ca9f9", x"060dedc9"),
	(x"88e10000", x"9ed20000", x"18d9c480", x"58660000", x"30c0573a", x"79b655db", x"01ec9988", x"34fbc344", x"0bf40000", x"f56c0001", x"42c13580", x"e2c30000", x"72203be1", x"48a08ee7", x"b2560bd4", x"886a5a33"),
	(x"bd480000", x"c51a0000", x"8d68ca00", x"66600000", x"578744be", x"c830d45b", x"7e79d306", x"13a978eb", x"c54f0000", x"e7270001", x"a2643100", x"8f0b0000", x"837d6dcd", x"4f737c98", x"7249578f", x"b6c637b6"),
	(x"715c0000", x"60790000", x"d7d1cd80", x"5d300000", x"1c575741", x"4fabe043", x"173a9bc7", x"d9f3ff15", x"44d10000", x"0b700001", x"c4563380", x"1af80000", x"ded445cf", x"07874024", x"9413f5a2", x"38a1804c"),
	(x"3cd60000", x"294d0000", x"eb5ac880", x"f3930000", x"0a2e6cbc", x"80c4e8e7", x"9823712b", x"9dcecf11", x"88c50000", x"ae130001", x"9eef3400", x"21a80000", x"95045630", x"801c743c", x"fd50bd63", x"f2fb07b2"),
	(x"f0c20000", x"8c2e0000", x"b1e3cf00", x"c8c30000", x"41fe7f43", x"075fdcff", x"f16039ea", x"579448ef", x"095b0000", x"42440001", x"f8dd3680", x"b45b0000", x"c8ad7e32", x"c8e84880", x"1b0a1f4e", x"7c9cb048"),
	(x"c7c40000", x"60ce0000", x"9e4ec280", x"a05d0000", x"9c342914", x"36919b18", x"27a967fe", x"8430193b", x"bd6c0000", x"f5db0001", x"0b5e3a80", x"1fae0000", x"f24345b4", x"319af5bc", x"82c5f7ed", x"d5a9bc1d"),
	(x"0bd00000", x"c5ad0000", x"c4f7c500", x"9b0d0000", x"d7e43aeb", x"b10aaf00", x"4eea2f3f", x"4e6a9ec5", x"3cf20000", x"198c0001", x"6d6c3800", x"8a5d0000", x"afea6db6", x"796ec900", x"649f55c0", x"5bce0be7"),
	(x"465a0000", x"8c990000", x"f87cc000", x"35ae0000", x"c19d0116", x"7e65a7a4", x"c1f3c5d3", x"0a57aec1", x"f0e60000", x"bcef0001", x"37d53f80", x"b10d0000", x"e43a7e49", x"fef5fd18", x"0ddc1d01", x"91948c19"),
	(x"8a4e0000", x"29fa0000", x"a2c5c780", x"0efe0000", x"8a4d12e9", x"f9fe93bc", x"a8b08d12", x"c00d293f", x"71780000", x"50b80001", x"51e73d00", x"24fe0000", x"b993564b", x"b601c1a4", x"eb86bf2c", x"1ff33be3"),
	(x"bfe70000", x"72320000", x"3774c900", x"30f80000", x"ed0a016d", x"4878123c", x"d725c79c", x"e75f9290", x"bfc30000", x"42f30001", x"b1423980", x"49360000", x"48ce0067", x"b1d233db", x"2b99e377", x"215f5666"),
	(x"73f30000", x"d7510000", x"6dcdce80", x"0ba80000", x"a6da1292", x"cfe32624", x"be668f5d", x"2d05156e", x"3e5d0000", x"aea40001", x"d7703b00", x"dcc50000", x"15672865", x"f9260f67", x"cdc3415a", x"af38e19c"),
	(x"3e790000", x"9e650000", x"5146cb80", x"a50b0000", x"b0a3296f", x"008c2e80", x"317f65b1", x"6938256a", x"f2490000", x"0bc70001", x"8dc93c80", x"e7950000", x"5eb73b9a", x"7ebd3b7f", x"a480099b", x"65626662"),
	(x"f26d0000", x"3b060000", x"0bffcc00", x"9e5b0000", x"fb733a90", x"87171a98", x"583c2d70", x"a362a294", x"73d70000", x"e7900001", x"ebfb3e00", x"72660000", x"031e1398", x"364907c3", x"42daabb6", x"eb05d198"),
	(x"69230000", x"cc400000", x"61a9d200", x"f5860000", x"7c3c5dad", x"a96b0dc9", x"7087b49a", x"e1228bb6", x"d9ae0000", x"8ec00001", x"75803380", x"aeb70000", x"d5b72f80", x"3b9bd3b1", x"16b65b07", x"da9a94a3"),
	(x"a5370000", x"69230000", x"3b10d580", x"ced60000", x"37ec4e52", x"2ef039d1", x"19c4fc5b", x"2b780c48", x"58300000", x"62970001", x"13b23100", x"3b440000", x"881e0782", x"736fef0d", x"f0ecf92a", x"54fd2359"),
	(x"e8bd0000", x"20170000", x"079bd080", x"60750000", x"219575af", x"e19f3175", x"96dd16b7", x"6f453c4c", x"94240000", x"c7f40001", x"490b3680", x"00140000", x"c3ce147d", x"f4f4db15", x"99afb1eb", x"9ea7a4a7"),
	(x"24a90000", x"85740000", x"5d22d700", x"5b250000", x"6a456650", x"6604056d", x"ff9e5e76", x"a51fbbb2", x"15ba0000", x"2ba30001", x"2f393400", x"95e70000", x"9e673c7f", x"bc00e7a9", x"7ff513c6", x"10c0135d"),
	(x"11000000", x"debc0000", x"c893d980", x"65230000", x"0d0275d4", x"d78284ed", x"800b14f8", x"824d001d", x"db010000", x"39e80001", x"cf9c3080", x"f82f0000", x"6f3a6a53", x"bbd315d6", x"bfea4f9d", x"2e6c7ed8"),
	(x"dd140000", x"7bdf0000", x"922ade00", x"5e730000", x"46d2662b", x"5019b0f5", x"e9485c39", x"481787e3", x"5a9f0000", x"d5bf0001", x"a9ae3200", x"6ddc0000", x"32934251", x"f327296a", x"59b0edb0", x"a00bc922"),
	(x"909e0000", x"32eb0000", x"aea1db00", x"f0d00000", x"50ab5dd6", x"9f76b851", x"6651b6d5", x"0c2ab7e7", x"968b0000", x"70dc0001", x"f3173580", x"568c0000", x"794351ae", x"74bc1d72", x"30f3a571", x"6a514edc"),
	(x"5c8a0000", x"97880000", x"f418dc80", x"cb800000", x"1b7b4e29", x"18ed8c49", x"0f12fe14", x"c6703019", x"17150000", x"9c8b0001", x"95253700", x"c37f0000", x"24ea79ac", x"3c4821ce", x"d6a9075c", x"e436f926"),
	(x"6b8c0000", x"7b680000", x"dbb5d100", x"a31e0000", x"c6b1187e", x"2923cbae", x"d9dba000", x"15d461cd", x"a3220000", x"2b140001", x"66a63b00", x"688a0000", x"1e04422a", x"c53a9cf2", x"4f66efff", x"4d03f573"),
	(x"a7980000", x"de0b0000", x"810cd680", x"984e0000", x"8d610b81", x"aeb8ffb6", x"b098e8c1", x"df8ee633", x"22bc0000", x"c7430001", x"00943980", x"fd790000", x"43ad6a28", x"8dcea04e", x"a93c4dd2", x"c3644289"),
	(x"ea120000", x"973f0000", x"bd87d380", x"36ed0000", x"9b18307c", x"61d7f712", x"3f81022d", x"9bb3d637", x"eea80000", x"62200001", x"5a2d3e00", x"c6290000", x"087d79d7", x"0a559456", x"c07f0513", x"093ec577"),
	(x"26060000", x"325c0000", x"e73ed400", x"0dbd0000", x"d0c82383", x"e64cc30a", x"56c24aec", x"51e951c9", x"6f360000", x"8e770001", x"3c1f3c80", x"53da0000", x"55d451d5", x"42a1a8ea", x"2625a73e", x"8759728d"),
	(x"13af0000", x"69940000", x"728fda80", x"33bb0000", x"b78f3007", x"57ca428a", x"29570062", x"76bbea66", x"a18d0000", x"9c3c0001", x"dcba3800", x"3e120000", x"a48907f9", x"45725a95", x"e63afb65", x"b9f51f08"),
	(x"dfbb0000", x"ccf70000", x"2836dd00", x"08eb0000", x"fc5f23f8", x"d0517692", x"401448a3", x"bce16d98", x"20130000", x"706b0001", x"ba883a80", x"abe10000", x"f9202ffb", x"0d866629", x"00605948", x"3792a8f2"),
	(x"92310000", x"85c30000", x"14bdd800", x"a6480000", x"ea261805", x"1f3e7e36", x"cf0da24f", x"f8dc5d9c", x"ec070000", x"d5080001", x"e0313d00", x"90b10000", x"b2f03c04", x"8a1d5231", x"69231189", x"fdc82f0c"),
	(x"5e250000", x"20a00000", x"4e04df80", x"9d180000", x"a1f60bfa", x"98a54a2e", x"a64eea8e", x"3286da62", x"6d990000", x"395f0001", x"86033f80", x"05420000", x"ef591406", x"c2e96e8d", x"8f79b3a4", x"73af98f6"),
	(x"75e60000", x"95660001", x"307b2000", x"adf40000", x"8f321eea", x"24298307", x"e8c49cf9", x"4b7eec55", x"aec30000", x"9c4f0001", x"79d1e000", x"2c150000", x"45cc75b3", x"6650b736", x"ab92f78f", x"a312567b"),
	(x"b9f20000", x"30050001", x"6ac22780", x"96a40000", x"c4e20d15", x"a3b2b71f", x"8187d438", x"81246bab", x"2f5d0000", x"70180001", x"1fe3e280", x"b9e60000", x"18655db1", x"2ea48b8a", x"4dc855a2", x"2d75e181"),
	(x"f4780000", x"79310001", x"56492280", x"38070000", x"d29b36e8", x"6cddbfbb", x"0e9e3ed4", x"c5195baf", x"e3490000", x"d57b0001", x"455ae500", x"82b60000", x"53b54e4e", x"a93fbf92", x"248b1d63", x"e72f667f"),
	(x"386c0000", x"dc520001", x"0cf02500", x"03570000", x"994b2517", x"eb468ba3", x"67dd7615", x"0f43dc51", x"62d70000", x"392c0001", x"2368e780", x"17450000", x"0e1c664c", x"e1cb832e", x"c2d1bf4e", x"6948d185"),
	(x"0dc50000", x"879a0001", x"99412b80", x"3d510000", x"fe0c3693", x"5ac00a23", x"18483c9b", x"281167fe", x"ac6c0000", x"2b670001", x"c3cde300", x"7a8d0000", x"ff413060", x"e6187151", x"02cee315", x"57e4bc00"),
	(x"c1d10000", x"22f90001", x"c3f82c00", x"06010000", x"b5dc256c", x"dd5b3e3b", x"710b745a", x"e24be000", x"2df20000", x"c7300001", x"a5ffe180", x"ef7e0000", x"a2e81862", x"aeec4ded", x"e4944138", x"d9830bfa"),
	(x"8c5b0000", x"6bcd0001", x"ff732900", x"a8a20000", x"a3a51e91", x"1234369f", x"fe129eb6", x"a676d004", x"e1e60000", x"62530001", x"ff46e600", x"d42e0000", x"e9380b9d", x"297779f5", x"8dd709f9", x"13d98c04"),
	(x"404f0000", x"ceae0001", x"a5ca2e80", x"93f20000", x"e8750d6e", x"95af0287", x"9751d677", x"6c2c57fa", x"60780000", x"8e040001", x"9974e480", x"41dd0000", x"b491239f", x"61834549", x"6b8dabd4", x"9dbe3bfe"),
	(x"77490000", x"224e0001", x"8a672300", x"fb6c0000", x"35bf5b39", x"a4614560", x"41988863", x"bf88062e", x"d44f0000", x"399b0001", x"6af7e880", x"ea280000", x"8e7f1819", x"98f1f875", x"f2424377", x"348b37ab"),
	(x"bb5d0000", x"872d0001", x"d0de2480", x"c03c0000", x"7e6f48c6", x"23fa7178", x"28dbc0a2", x"75d281d0", x"55d10000", x"d5cc0001", x"0cc5ea00", x"7fdb0000", x"d3d6301b", x"d005c4c9", x"1418e15a", x"baec8051"),
	(x"f6d70000", x"ce190001", x"ec552180", x"6e9f0000", x"6816733b", x"ec9579dc", x"a7c22a4e", x"31efb1d4", x"99c50000", x"70af0001", x"567ced80", x"448b0000", x"980623e4", x"579ef0d1", x"7d5ba99b", x"70b607af"),
	(x"3ac30000", x"6b7a0001", x"b6ec2600", x"55cf0000", x"23c660c4", x"6b0e4dc4", x"ce81628f", x"fbb5362a", x"185b0000", x"9cf80001", x"304eef00", x"d1780000", x"c5af0be6", x"1f6acc6d", x"9b010bb6", x"fed1b055"),
	(x"0f6a0000", x"30b20001", x"235d2880", x"6bc90000", x"44817340", x"da88cc44", x"b1142801", x"dce78d85", x"d6e00000", x"8eb30001", x"d0ebeb80", x"bcb00000", x"34f25dca", x"18b93e12", x"5b1e57ed", x"c07dddd0"),
	(x"c37e0000", x"95d10001", x"79e42f00", x"50990000", x"0f5160bf", x"5d13f85c", x"d85760c0", x"16bd0a7b", x"577e0000", x"62e40001", x"b6d9e900", x"29430000", x"695b75c8", x"504d02ae", x"bd44f5c0", x"4e1a6a2a"),
	(x"8ef40000", x"dce50001", x"456f2a00", x"fe3a0000", x"19285b42", x"927cf0f8", x"574e8a2c", x"52803a7f", x"9b6a0000", x"c7870001", x"ec60ee80", x"12130000", x"228b6637", x"d7d636b6", x"d407bd01", x"8440edd4"),
	(x"42e00000", x"79860001", x"1fd62d80", x"c56a0000", x"52f848bd", x"15e7c4e0", x"3e0dc2ed", x"98dabd81", x"1af40000", x"2bd00001", x"8a52ec00", x"87e00000", x"7f224e35", x"9f220a0a", x"325d1f2c", x"0a275a2e"),
	(x"d9ae0000", x"8ec00001", x"75803380", x"aeb70000", x"d5b72f80", x"3b9bd3b1", x"16b65b07", x"da9a94a3", x"b08d0000", x"42800001", x"1429e180", x"5b310000", x"a98b722d", x"92f0de78", x"6631ef9d", x"3bb81f15"),
	(x"15ba0000", x"2ba30001", x"2f393400", x"95e70000", x"9e673c7f", x"bc00e7a9", x"7ff513c6", x"10c0135d", x"31130000", x"aed70001", x"721be300", x"cec20000", x"f4225a2f", x"da04e2c4", x"806b4db0", x"b5dfa8ef"),
	(x"58300000", x"62970001", x"13b23100", x"3b440000", x"881e0782", x"736fef0d", x"f0ecf92a", x"54fd2359", x"fd070000", x"0bb40001", x"28a2e480", x"f5920000", x"bff249d0", x"5d9fd6dc", x"e9280571", x"7f852f11"),
	(x"94240000", x"c7f40001", x"490b3680", x"00140000", x"c3ce147d", x"f4f4db15", x"99afb1eb", x"9ea7a4a7", x"7c990000", x"e7e30001", x"4e90e600", x"60610000", x"e25b61d2", x"156bea60", x"0f72a75c", x"f1e298eb"),
	(x"a18d0000", x"9c3c0001", x"dcba3800", x"3e120000", x"a48907f9", x"45725a95", x"e63afb65", x"b9f51f08", x"b2220000", x"f5a80001", x"ae35e280", x"0da90000", x"130637fe", x"12b8181f", x"cf6dfb07", x"cf4ef56e"),
	(x"6d990000", x"395f0001", x"86033f80", x"05420000", x"ef591406", x"c2e96e8d", x"8f79b3a4", x"73af98f6", x"33bc0000", x"19ff0001", x"c807e000", x"985a0000", x"4eaf1ffc", x"5a4c24a3", x"2937592a", x"41294294"),
	(x"20130000", x"706b0001", x"ba883a80", x"abe10000", x"f9202ffb", x"0d866629", x"00605948", x"3792a8f2", x"ffa80000", x"bc9c0001", x"92bee780", x"a30a0000", x"057f0c03", x"ddd710bb", x"407411eb", x"8b73c56a"),
	(x"ec070000", x"d5080001", x"e0313d00", x"90b10000", x"b2f03c04", x"8a1d5231", x"69231189", x"fdc82f0c", x"7e360000", x"50cb0001", x"f48ce500", x"36f90000", x"58d62401", x"95232c07", x"a62eb3c6", x"05147290"),
	(x"db010000", x"39e80001", x"cf9c3080", x"f82f0000", x"6f3a6a53", x"bbd315d6", x"bfea4f9d", x"2e6c7ed8", x"ca010000", x"e7540001", x"070fe900", x"9d0c0000", x"62381f87", x"6c51913b", x"3fe15b65", x"ac217ec5"),
	(x"17150000", x"9c8b0001", x"95253700", x"c37f0000", x"24ea79ac", x"3c4821ce", x"d6a9075c", x"e436f926", x"4b9f0000", x"0b030001", x"613deb80", x"08ff0000", x"3f913785", x"24a5ad87", x"d9bbf948", x"2246c93f"),
	(x"5a9f0000", x"d5bf0001", x"a9ae3200", x"6ddc0000", x"32934251", x"f327296a", x"59b0edb0", x"a00bc922", x"878b0000", x"ae600001", x"3b84ec00", x"33af0000", x"7441247a", x"a33e999f", x"b0f8b189", x"e81c4ec1"),
	(x"968b0000", x"70dc0001", x"f3173580", x"568c0000", x"794351ae", x"74bc1d72", x"30f3a571", x"6a514edc", x"06150000", x"42370001", x"5db6ee80", x"a65c0000", x"29e80c78", x"ebcaa523", x"56a213a4", x"667bf93b"),
	(x"a3220000", x"2b140001", x"66a63b00", x"688a0000", x"1e04422a", x"c53a9cf2", x"4f66efff", x"4d03f573", x"c8ae0000", x"507c0001", x"bd13ea00", x"cb940000", x"d8b55a54", x"ec19575c", x"96bd4fff", x"58d794be"),
	(x"6f360000", x"8e770001", x"3c1f3c80", x"53da0000", x"55d451d5", x"42a1a8ea", x"2625a73e", x"8759728d", x"49300000", x"bc2b0001", x"db21e880", x"5e670000", x"851c7256", x"a4ed6be0", x"70e7edd2", x"d6b02344"),
	(x"22bc0000", x"c7430001", x"00943980", x"fd790000", x"43ad6a28", x"8dcea04e", x"a93c4dd2", x"c3644289", x"85240000", x"19480001", x"8198ef00", x"65370000", x"cecc61a9", x"23765ff8", x"19a4a513", x"1ceaa4ba"),
	(x"eea80000", x"62200001", x"5a2d3e00", x"c6290000", x"087d79d7", x"0a559456", x"c07f0513", x"093ec577", x"04ba0000", x"f51f0001", x"e7aaed80", x"f0c40000", x"936549ab", x"6b826344", x"fffe073e", x"928d1340"),
	(x"6ba80000", x"4ba90001", x"5d832180", x"dad00000", x"63751974", x"d089ea49", x"256784eb", x"d3d4a53b", x"1cc50000", x"59260001", x"51d2f200", x"58720000", x"f30e4347", x"8d428ece", x"98432863", x"aa5c67e3"),
	(x"a7bc0000", x"eeca0001", x"073a2600", x"e1800000", x"28a50a8b", x"5712de51", x"4c24cc2a", x"198e22c5", x"9d5b0000", x"b5710001", x"37e0f080", x"cd810000", x"aea76b45", x"c5b6b272", x"7e198a4e", x"243bd019"),
	(x"ea360000", x"a7fe0001", x"3bb12300", x"4f230000", x"3edc3176", x"987dd6f5", x"c33d26c6", x"5db312c1", x"514f0000", x"10120001", x"6d59f700", x"f6d10000", x"e57778ba", x"422d866a", x"175ac28f", x"ee6157e7"),
	(x"26220000", x"029d0001", x"61082480", x"74730000", x"750c2289", x"1fe6e2ed", x"aa7e6e07", x"97e9953f", x"d0d10000", x"fc450001", x"0b6bf580", x"63220000", x"b8de50b8", x"0ad9bad6", x"f10060a2", x"6006e01d"),
	(x"138b0000", x"59550001", x"f4b92a00", x"4a750000", x"124b310d", x"ae60636d", x"d5eb2489", x"b0bb2e90", x"1e6a0000", x"ee0e0001", x"ebcef100", x"0eea0000", x"49830694", x"0d0a48a9", x"311f3cf9", x"5eaa8d98"),
	(x"df9f0000", x"fc360001", x"ae002d80", x"71250000", x"599b22f2", x"29fb5775", x"bca86c48", x"7ae1a96e", x"9ff40000", x"02590001", x"8dfcf380", x"9b190000", x"142a2e96", x"45fe7415", x"d7459ed4", x"d0cd3a62"),
	(x"92150000", x"b5020001", x"928b2880", x"df860000", x"4fe2190f", x"e6945fd1", x"33b186a4", x"3edc996a", x"53e00000", x"a73a0001", x"d745f400", x"a0490000", x"5ffa3d69", x"c265400d", x"be06d615", x"1a97bd9c"),
	(x"5e010000", x"10610001", x"c8322f00", x"e4d60000", x"04320af0", x"610f6bc9", x"5af2ce65", x"f4861e94", x"d27e0000", x"4b6d0001", x"b177f680", x"35ba0000", x"0253156b", x"8a917cb1", x"585c7438", x"94f00a66"),
	(x"69070000", x"fc810001", x"e79f2280", x"8c480000", x"d9f85ca7", x"50c12c2e", x"8c3b9071", x"27224f40", x"66490000", x"fcf20001", x"42f4fa80", x"9e4f0000", x"38bd2eed", x"73e3c18d", x"c1939c9b", x"3dc50633"),
	(x"a5130000", x"59e20001", x"bd262500", x"b7180000", x"92284f58", x"d75a1836", x"e578d8b0", x"ed78c8be", x"e7d70000", x"10a50001", x"24c6f800", x"0bbc0000", x"651406ef", x"3b17fd31", x"27c93eb6", x"b3a2b1c9"),
	(x"e8990000", x"10d60001", x"81ad2000", x"19bb0000", x"845174a5", x"18351092", x"6a61325c", x"a945f8ba", x"2bc30000", x"b5c60001", x"7e7fff80", x"30ec0000", x"2ec41510", x"bc8cc929", x"4e8a7677", x"79f83637"),
	(x"248d0000", x"b5b50001", x"db142780", x"22eb0000", x"cf81675a", x"9fae248a", x"03227a9d", x"631f7f44", x"aa5d0000", x"59910001", x"184dfd00", x"a51f0000", x"736d3d12", x"f478f595", x"a8d0d45a", x"f79f81cd"),
	(x"11240000", x"ee7d0001", x"4ea52900", x"1ced0000", x"a8c674de", x"2e28a50a", x"7cb73013", x"444dc4eb", x"64e60000", x"4bda0001", x"f8e8f980", x"c8d70000", x"82306b3e", x"f3ab07ea", x"68cf8801", x"c933ec48"),
	(x"dd300000", x"4b1e0001", x"141c2e80", x"27bd0000", x"e3166721", x"a9b39112", x"15f478d2", x"8e174315", x"e5780000", x"a78d0001", x"9edafb00", x"5d240000", x"df99433c", x"bb5f3b56", x"8e952a2c", x"47545bb2"),
	(x"90ba0000", x"022a0001", x"28972b80", x"891e0000", x"f56f5cdc", x"66dc99b6", x"9aed923e", x"ca2a7311", x"296c0000", x"02ee0001", x"c463fc80", x"66740000", x"944950c3", x"3cc40f4e", x"e7d662ed", x"8d0edc4c"),
	(x"5cae0000", x"a7490001", x"722e2c00", x"b24e0000", x"bebf4f23", x"e147adae", x"f3aedaff", x"0070f4ef", x"a8f20000", x"eeb90001", x"a251fe00", x"f3870000", x"c9e078c1", x"743033f2", x"018cc0c0", x"03696bb6"),
	(x"c7e00000", x"500f0001", x"18783200", x"d9930000", x"39f0281e", x"cf3bbaff", x"db154315", x"4230ddcd", x"028b0000", x"87e90001", x"3c2af380", x"2f560000", x"1f4944d9", x"79e2e780", x"55e03071", x"32f62e8d"),
	(x"0bf40000", x"f56c0001", x"42c13580", x"e2c30000", x"72203be1", x"48a08ee7", x"b2560bd4", x"886a5a33", x"83150000", x"6bbe0001", x"5a18f100", x"baa50000", x"42e06cdb", x"3116db3c", x"b3ba925c", x"bc919977"),
	(x"467e0000", x"bc580001", x"7e4a3080", x"4c600000", x"6459001c", x"87cf8643", x"3d4fe138", x"cc576a37", x"4f010000", x"cedd0001", x"00a1f680", x"81f50000", x"09307f24", x"b68def24", x"daf9da9d", x"76cb1e89"),
	(x"8a6a0000", x"193b0001", x"24f33700", x"77300000", x"2f8913e3", x"0054b25b", x"540ca9f9", x"060dedc9", x"ce9f0000", x"228a0001", x"6693f400", x"14060000", x"54995726", x"fe79d398", x"3ca378b0", x"f8aca973"),
	(x"bfc30000", x"42f30001", x"b1423980", x"49360000", x"48ce0067", x"b1d233db", x"2b99e377", x"215f5666", x"00240000", x"30c10001", x"8636f080", x"79ce0000", x"a5c4010a", x"f9aa21e7", x"fcbc24eb", x"c600c4f6"),
	(x"73d70000", x"e7900001", x"ebfb3e00", x"72660000", x"031e1398", x"364907c3", x"42daabb6", x"eb05d198", x"81ba0000", x"dc960001", x"e004f200", x"ec3d0000", x"f86d2908", x"b15e1d5b", x"1ae686c6", x"4867730c"),
	(x"3e5d0000", x"aea40001", x"d7703b00", x"dcc50000", x"15672865", x"f9260f67", x"cdc3415a", x"af38e19c", x"4dae0000", x"79f50001", x"babdf580", x"d76d0000", x"b3bd3af7", x"36c52943", x"73a5ce07", x"823df4f2"),
	(x"f2490000", x"0bc70001", x"8dc93c80", x"e7950000", x"5eb73b9a", x"7ebd3b7f", x"a480099b", x"65626662", x"cc300000", x"95a20001", x"dc8ff700", x"429e0000", x"ee1412f5", x"7e3115ff", x"95ff6c2a", x"0c5a4308"),
	(x"c54f0000", x"e7270001", x"a2643100", x"8f0b0000", x"837d6dcd", x"4f737c98", x"7249578f", x"b6c637b6", x"78070000", x"223d0001", x"2f0cfb00", x"e96b0000", x"d4fa2973", x"8743a8c3", x"0c308489", x"a56f4f5d"),
	(x"095b0000", x"42440001", x"f8dd3680", x"b45b0000", x"c8ad7e32", x"c8e84880", x"1b0a1f4e", x"7c9cb048", x"f9990000", x"ce6a0001", x"493ef980", x"7c980000", x"89530171", x"cfb7947f", x"ea6a26a4", x"2b08f8a7"),
	(x"44d10000", x"0b700001", x"c4563380", x"1af80000", x"ded445cf", x"07874024", x"9413f5a2", x"38a1804c", x"358d0000", x"6b090001", x"1387fe00", x"47c80000", x"c283128e", x"482ca067", x"83296e65", x"e1527f59"),
	(x"88c50000", x"ae130001", x"9eef3400", x"21a80000", x"95045630", x"801c743c", x"fd50bd63", x"f2fb07b2", x"b4130000", x"875e0001", x"75b5fc80", x"d23b0000", x"9f2a3a8c", x"00d89cdb", x"6573cc48", x"6f35c8a3"),
	(x"bd6c0000", x"f5db0001", x"0b5e3a80", x"1fae0000", x"f24345b4", x"319af5bc", x"82c5f7ed", x"d5a9bc1d", x"7aa80000", x"95150001", x"9510f800", x"bff30000", x"6e776ca0", x"070b6ea4", x"a56c9013", x"5199a526"),
	(x"71780000", x"50b80001", x"51e73d00", x"24fe0000", x"b993564b", x"b601c1a4", x"eb86bf2c", x"1ff33be3", x"fb360000", x"79420001", x"f322fa80", x"2a000000", x"33de44a2", x"4fff5218", x"4336323e", x"dffe12dc"),
	(x"3cf20000", x"198c0001", x"6d6c3800", x"8a5d0000", x"afea6db6", x"796ec900", x"649f55c0", x"5bce0be7", x"37220000", x"dc210001", x"a99bfd00", x"11500000", x"780e575d", x"c8646600", x"2a757aff", x"15a49522"),
	(x"f0e60000", x"bcef0001", x"37d53f80", x"b10d0000", x"e43a7e49", x"fef5fd18", x"0ddc1d01", x"91948c19", x"b6bc0000", x"30760001", x"cfa9ff80", x"84a30000", x"25a77f5f", x"80905abc", x"cc2fd8d2", x"9bc322d8")
    ),(
	(x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000"),
	(x"58430000", x"807e0000", x"78330001", x"c66b3800", x"e7375cdc", x"79ad3fdd", x"ac73fe6f", x"3a4479b1", x"1d5a0000", x"2b720000", x"488d0000", x"af611800", x"25cb2ec5", x"c879bfd0", x"81a20429", x"1e7536a6"),
	(x"1d5a0000", x"2b720000", x"488d0000", x"af611800", x"25cb2ec5", x"c879bfd0", x"81a20429", x"1e7536a6", x"45190000", x"ab0c0000", x"30be0001", x"690a2000", x"c2fc7219", x"b1d4800d", x"2dd1fa46", x"24314f17"),
	(x"45190000", x"ab0c0000", x"30be0001", x"690a2000", x"c2fc7219", x"b1d4800d", x"2dd1fa46", x"24314f17", x"58430000", x"807e0000", x"78330001", x"c66b3800", x"e7375cdc", x"79ad3fdd", x"ac73fe6f", x"3a4479b1"),
	(x"a53b0000", x"14260000", x"4e30001e", x"7cae0000", x"8f9e0dd5", x"78dfaa3d", x"f73168d8", x"0b1b4946", x"07ed0000", x"b2500000", x"8774000a", x"970d0000", x"437223ae", x"48c76ea4", x"f4786222", x"9075b1ce"),
	(x"fd780000", x"94580000", x"3603001f", x"bac53800", x"68a95109", x"017295e0", x"5b4296b7", x"315f30f7", x"1ab70000", x"99220000", x"cff9000a", x"386c1800", x"66b90d6b", x"80bed174", x"75da660b", x"8e008768"),
	(x"b8610000", x"3f540000", x"06bd001e", x"d3cf1800", x"aa552310", x"b0a615ed", x"76936cf1", x"156e7fe0", x"42f40000", x"195c0000", x"b7ca000b", x"fe072000", x"818e51b7", x"f913eea9", x"d9a99864", x"b444fed9"),
	(x"e0220000", x"bf2a0000", x"7e8e001f", x"15a42000", x"4d627fcc", x"c90b2a30", x"dae0929e", x"2f2a0651", x"5fae0000", x"322e0000", x"ff47000b", x"51663800", x"a4457f72", x"316a5179", x"580b9c4d", x"aa31c87f"),
	(x"07ed0000", x"b2500000", x"8774000a", x"970d0000", x"437223ae", x"48c76ea4", x"f4786222", x"9075b1ce", x"a2d60000", x"a6760000", x"c9440014", x"eba30000", x"ccec2e7b", x"3018c499", x"03490afa", x"9b6ef888"),
	(x"5fae0000", x"322e0000", x"ff47000b", x"51663800", x"a4457f72", x"316a5179", x"580b9c4d", x"aa31c87f", x"bf8c0000", x"8d040000", x"81c90014", x"44c21800", x"e92700be", x"f8617b49", x"82eb0ed3", x"851bce2e"),
	(x"1ab70000", x"99220000", x"cff9000a", x"386c1800", x"66b90d6b", x"80bed174", x"75da660b", x"8e008768", x"e7cf0000", x"0d7a0000", x"f9fa0015", x"82a92000", x"0e105c62", x"81cc4494", x"2e98f0bc", x"bf5fb79f"),
	(x"42f40000", x"195c0000", x"b7ca000b", x"fe072000", x"818e51b7", x"f913eea9", x"d9a99864", x"b444fed9", x"fa950000", x"26080000", x"b1770015", x"2dc83800", x"2bdb72a7", x"49b5fb44", x"af3af495", x"a12a8139"),
	(x"a2d60000", x"a6760000", x"c9440014", x"eba30000", x"ccec2e7b", x"3018c499", x"03490afa", x"9b6ef888", x"a53b0000", x"14260000", x"4e30001e", x"7cae0000", x"8f9e0dd5", x"78dfaa3d", x"f73168d8", x"0b1b4946"),
	(x"fa950000", x"26080000", x"b1770015", x"2dc83800", x"2bdb72a7", x"49b5fb44", x"af3af495", x"a12a8139", x"b8610000", x"3f540000", x"06bd001e", x"d3cf1800", x"aa552310", x"b0a615ed", x"76936cf1", x"156e7fe0"),
	(x"bf8c0000", x"8d040000", x"81c90014", x"44c21800", x"e92700be", x"f8617b49", x"82eb0ed3", x"851bce2e", x"e0220000", x"bf2a0000", x"7e8e001f", x"15a42000", x"4d627fcc", x"c90b2a30", x"dae0929e", x"2f2a0651"),
	(x"e7cf0000", x"0d7a0000", x"f9fa0015", x"82a92000", x"0e105c62", x"81cc4494", x"2e98f0bc", x"bf5fb79f", x"fd780000", x"94580000", x"3603001f", x"bac53800", x"68a95109", x"017295e0", x"5b4296b7", x"315f30f7"),
	(x"88980000", x"1f940000", x"7fcf002e", x"fb4e0000", x"f158079a", x"61ae9167", x"a895706c", x"e6107494", x"0bc20000", x"db630000", x"7e88000c", x"15860000", x"91fd48f3", x"7581bb43", x"f460449e", x"d8b61463"),
	(x"d0db0000", x"9fea0000", x"07fc002f", x"3d253800", x"166f5b46", x"1803aeba", x"04e68e03", x"dc540d25", x"16980000", x"f0110000", x"3605000c", x"bae71800", x"b4366636", x"bdf80493", x"75c240b7", x"c6c322c5"),
	(x"95c20000", x"34e60000", x"3742002e", x"542f1800", x"d493295f", x"a9d72eb7", x"29377445", x"f8654232", x"4edb0000", x"706f0000", x"4e36000d", x"7c8c2000", x"53013aea", x"c4553b4e", x"d9b1bed8", x"fc875b74"),
	(x"cd810000", x"b4980000", x"4f71002f", x"92442000", x"33a47583", x"d07a116a", x"85448a2a", x"c2213b83", x"53810000", x"5b1d0000", x"06bb000d", x"d3ed3800", x"76ca142f", x"0c2c849e", x"5813baf1", x"e2f26dd2"),
	(x"2da30000", x"0bb20000", x"31ff0030", x"87e00000", x"7ec60a4f", x"19713b5a", x"5fa418b4", x"ed0b3dd2", x"0c2f0000", x"69330000", x"f9fc0006", x"828b0000", x"d28f6b5d", x"3d46d5e7", x"001826bc", x"48c3a5ad"),
	(x"75e00000", x"8bcc0000", x"49cc0031", x"418b3800", x"99f15693", x"60dc0487", x"f3d7e6db", x"d74f4463", x"11750000", x"42410000", x"b1710006", x"2dea1800", x"f7444598", x"f53f6a37", x"81ba2295", x"56b6930b"),
	(x"30f90000", x"20c00000", x"79720030", x"28811800", x"5b0d248a", x"d108848a", x"de061c9d", x"f37e0b74", x"49360000", x"c23f0000", x"c9420007", x"eb812000", x"10731944", x"8c9255ea", x"2dc9dcfa", x"6cf2eaba"),
	(x"68ba0000", x"a0be0000", x"01410031", x"eeea2000", x"bc3a7856", x"a8a5bb57", x"7275e2f2", x"c93a72c5", x"546c0000", x"e94d0000", x"81cf0007", x"44e03800", x"35b83781", x"44ebea3a", x"ac6bd8d3", x"7287dc1c"),
	(x"8f750000", x"adc40000", x"f8bb0024", x"6c430000", x"b22a2434", x"2969ffc3", x"5ced124e", x"7665c55a", x"a9140000", x"7d150000", x"b7cc0018", x"fe250000", x"5d116688", x"45997fda", x"f7294e64", x"43d8eceb"),
	(x"d7360000", x"2dba0000", x"80880025", x"aa283800", x"551d78e8", x"50c4c01e", x"f09eec21", x"4c21bceb", x"b44e0000", x"56670000", x"ff410018", x"51441800", x"78da484d", x"8de0c00a", x"768b4a4d", x"5dadda4d"),
	(x"922f0000", x"86b60000", x"b0360024", x"c3221800", x"97e10af1", x"e1104013", x"dd4f1667", x"6810f3fc", x"ec0d0000", x"d6190000", x"87720019", x"972f2000", x"9fed1491", x"f44dffd7", x"daf8b422", x"67e9a3fc"),
	(x"ca6c0000", x"06c80000", x"c8050025", x"05492000", x"70d6562d", x"98bd7fce", x"713ce808", x"52548a4d", x"f1570000", x"fd6b0000", x"cfff0019", x"384e3800", x"ba263a54", x"3c344007", x"5b5ab00b", x"799c955a"),
	(x"2a4e0000", x"b9e20000", x"b68b003a", x"10ed0000", x"3db429e1", x"51b655fe", x"abdc7a96", x"7d7e8c1c", x"aef90000", x"cf450000", x"30b80012", x"69280000", x"1e634526", x"0d5e117e", x"03512c46", x"d3ad5d25"),
	(x"720d0000", x"399c0000", x"ceb8003b", x"d6863800", x"da83753d", x"281b6a23", x"07af84f9", x"473af5ad", x"b3a30000", x"e4370000", x"78350012", x"c6491800", x"3ba86be3", x"c527aeae", x"82f3286f", x"cdd86b83"),
	(x"37140000", x"92900000", x"fe06003a", x"bf8c1800", x"187f0724", x"99cfea2e", x"2a7e7ebf", x"630bbaba", x"ebe00000", x"64490000", x"00060013", x"00222000", x"dc9f373f", x"bc8a9173", x"2e80d600", x"f79c1232"),
	(x"6f570000", x"12ee0000", x"8635003b", x"79e72000", x"ff485bf8", x"e062d5f3", x"860d80d0", x"594fc30b", x"f6ba0000", x"4f3b0000", x"488b0013", x"af433800", x"f95419fa", x"74f32ea3", x"af22d229", x"e9e92494"),
	(x"0bc20000", x"db630000", x"7e88000c", x"15860000", x"91fd48f3", x"7581bb43", x"f460449e", x"d8b61463", x"835a0000", x"c4f70000", x"01470022", x"eec80000", x"60a54f69", x"142f2a24", x"5cf534f2", x"3ea660f7"),
	(x"53810000", x"5b1d0000", x"06bb000d", x"d3ed3800", x"76ca142f", x"0c2c849e", x"5813baf1", x"e2f26dd2", x"9e000000", x"ef850000", x"49ca0022", x"41a91800", x"456e61ac", x"dc5695f4", x"dd5730db", x"20d35651"),
	(x"16980000", x"f0110000", x"3605000c", x"bae71800", x"b4366636", x"bdf80493", x"75c240b7", x"c6c322c5", x"c6430000", x"6ffb0000", x"31f90023", x"87c22000", x"a2593d70", x"a5fbaa29", x"7124ceb4", x"1a972fe0"),
	(x"4edb0000", x"706f0000", x"4e36000d", x"7c8c2000", x"53013aea", x"c4553b4e", x"d9b1bed8", x"fc875b74", x"db190000", x"44890000", x"79740023", x"28a33800", x"879213b5", x"6d8215f9", x"f086ca9d", x"04e21946"),
	(x"aef90000", x"cf450000", x"30b80012", x"69280000", x"1e634526", x"0d5e117e", x"03512c46", x"d3ad5d25", x"84b70000", x"76a70000", x"86330028", x"79c50000", x"23d76cc7", x"5ce84480", x"a88d56d0", x"aed3d139"),
	(x"f6ba0000", x"4f3b0000", x"488b0013", x"af433800", x"f95419fa", x"74f32ea3", x"af22d229", x"e9e92494", x"99ed0000", x"5dd50000", x"cebe0028", x"d6a41800", x"061c4202", x"9491fb50", x"292f52f9", x"b0a6e79f"),
	(x"b3a30000", x"e4370000", x"78350012", x"c6491800", x"3ba86be3", x"c527aeae", x"82f3286f", x"cdd86b83", x"c1ae0000", x"ddab0000", x"b68d0029", x"10cf2000", x"e12b1ede", x"ed3cc48d", x"855cac96", x"8ae29e2e"),
	(x"ebe00000", x"64490000", x"00060013", x"00222000", x"dc9f373f", x"bc8a9173", x"2e80d600", x"f79c1232", x"dcf40000", x"f6d90000", x"fe000029", x"bfae3800", x"c4e0301b", x"25457b5d", x"04fea8bf", x"9497a888"),
	(x"0c2f0000", x"69330000", x"f9fc0006", x"828b0000", x"d28f6b5d", x"3d46d5e7", x"001826bc", x"48c3a5ad", x"218c0000", x"62810000", x"c8030036", x"056b0000", x"ac496112", x"2437eebd", x"5fbc3e08", x"a5c8987f"),
	(x"546c0000", x"e94d0000", x"81cf0007", x"44e03800", x"35b83781", x"44ebea3a", x"ac6bd8d3", x"7287dc1c", x"3cd60000", x"49f30000", x"808e0036", x"aa0a1800", x"89824fd7", x"ec4e516d", x"de1e3a21", x"bbbdaed9"),
	(x"11750000", x"42410000", x"b1710006", x"2dea1800", x"f7444598", x"f53f6a37", x"81ba2295", x"56b6930b", x"64950000", x"c98d0000", x"f8bd0037", x"6c612000", x"6eb5130b", x"95e36eb0", x"726dc44e", x"81f9d768"),
	(x"49360000", x"c23f0000", x"c9420007", x"eb812000", x"10731944", x"8c9255ea", x"2dc9dcfa", x"6cf2eaba", x"79cf0000", x"e2ff0000", x"b0300037", x"c3003800", x"4b7e3dce", x"5d9ad160", x"f3cfc067", x"9f8ce1ce"),
	(x"a9140000", x"7d150000", x"b7cc0018", x"fe250000", x"5d116688", x"45997fda", x"f7294e64", x"43d8eceb", x"26610000", x"d0d10000", x"4f77003c", x"92660000", x"ef3b42bc", x"6cf08019", x"abc45c2a", x"35bd29b1"),
	(x"f1570000", x"fd6b0000", x"cfff0019", x"384e3800", x"ba263a54", x"3c344007", x"5b5ab00b", x"799c955a", x"3b3b0000", x"fba30000", x"07fa003c", x"3d071800", x"caf06c79", x"a4893fc9", x"2a665803", x"2bc81f17"),
	(x"b44e0000", x"56670000", x"ff410018", x"51441800", x"78da484d", x"8de0c00a", x"768b4a4d", x"5dadda4d", x"63780000", x"7bdd0000", x"7fc9003d", x"fb6c2000", x"2dc730a5", x"dd240014", x"8615a66c", x"118c66a6"),
	(x"ec0d0000", x"d6190000", x"87720019", x"972f2000", x"9fed1491", x"f44dffd7", x"daf8b422", x"67e9a3fc", x"7e220000", x"50af0000", x"3744003d", x"540d3800", x"080c1e60", x"155dbfc4", x"07b7a245", x"0ff95000"),
	(x"835a0000", x"c4f70000", x"01470022", x"eec80000", x"60a54f69", x"142f2a24", x"5cf534f2", x"3ea660f7", x"88980000", x"1f940000", x"7fcf002e", x"fb4e0000", x"f158079a", x"61ae9167", x"a895706c", x"e6107494"),
	(x"db190000", x"44890000", x"79740023", x"28a33800", x"879213b5", x"6d8215f9", x"f086ca9d", x"04e21946", x"95c20000", x"34e60000", x"3742002e", x"542f1800", x"d493295f", x"a9d72eb7", x"29377445", x"f8654232"),
	(x"9e000000", x"ef850000", x"49ca0022", x"41a91800", x"456e61ac", x"dc5695f4", x"dd5730db", x"20d35651", x"cd810000", x"b4980000", x"4f71002f", x"92442000", x"33a47583", x"d07a116a", x"85448a2a", x"c2213b83"),
	(x"c6430000", x"6ffb0000", x"31f90023", x"87c22000", x"a2593d70", x"a5fbaa29", x"7124ceb4", x"1a972fe0", x"d0db0000", x"9fea0000", x"07fc002f", x"3d253800", x"166f5b46", x"1803aeba", x"04e68e03", x"dc540d25"),
	(x"26610000", x"d0d10000", x"4f77003c", x"92660000", x"ef3b42bc", x"6cf08019", x"abc45c2a", x"35bd29b1", x"8f750000", x"adc40000", x"f8bb0024", x"6c430000", x"b22a2434", x"2969ffc3", x"5ced124e", x"7665c55a"),
	(x"7e220000", x"50af0000", x"3744003d", x"540d3800", x"080c1e60", x"155dbfc4", x"07b7a245", x"0ff95000", x"922f0000", x"86b60000", x"b0360024", x"c3221800", x"97e10af1", x"e1104013", x"dd4f1667", x"6810f3fc"),
	(x"3b3b0000", x"fba30000", x"07fa003c", x"3d071800", x"caf06c79", x"a4893fc9", x"2a665803", x"2bc81f17", x"ca6c0000", x"06c80000", x"c8050025", x"05492000", x"70d6562d", x"98bd7fce", x"713ce808", x"52548a4d"),
	(x"63780000", x"7bdd0000", x"7fc9003d", x"fb6c2000", x"2dc730a5", x"dd240014", x"8615a66c", x"118c66a6", x"d7360000", x"2dba0000", x"80880025", x"aa283800", x"551d78e8", x"50c4c01e", x"f09eec21", x"4c21bceb"),
	(x"84b70000", x"76a70000", x"86330028", x"79c50000", x"23d76cc7", x"5ce84480", x"a88d56d0", x"aed3d139", x"2a4e0000", x"b9e20000", x"b68b003a", x"10ed0000", x"3db429e1", x"51b655fe", x"abdc7a96", x"7d7e8c1c"),
	(x"dcf40000", x"f6d90000", x"fe000029", x"bfae3800", x"c4e0301b", x"25457b5d", x"04fea8bf", x"9497a888", x"37140000", x"92900000", x"fe06003a", x"bf8c1800", x"187f0724", x"99cfea2e", x"2a7e7ebf", x"630bbaba"),
	(x"99ed0000", x"5dd50000", x"cebe0028", x"d6a41800", x"061c4202", x"9491fb50", x"292f52f9", x"b0a6e79f", x"6f570000", x"12ee0000", x"8635003b", x"79e72000", x"ff485bf8", x"e062d5f3", x"860d80d0", x"594fc30b"),
	(x"c1ae0000", x"ddab0000", x"b68d0029", x"10cf2000", x"e12b1ede", x"ed3cc48d", x"855cac96", x"8ae29e2e", x"720d0000", x"399c0000", x"ceb8003b", x"d6863800", x"da83753d", x"281b6a23", x"07af84f9", x"473af5ad"),
	(x"218c0000", x"62810000", x"c8030036", x"056b0000", x"ac496112", x"2437eebd", x"5fbc3e08", x"a5c8987f", x"2da30000", x"0bb20000", x"31ff0030", x"87e00000", x"7ec60a4f", x"19713b5a", x"5fa418b4", x"ed0b3dd2"),
	(x"79cf0000", x"e2ff0000", x"b0300037", x"c3003800", x"4b7e3dce", x"5d9ad160", x"f3cfc067", x"9f8ce1ce", x"30f90000", x"20c00000", x"79720030", x"28811800", x"5b0d248a", x"d108848a", x"de061c9d", x"f37e0b74"),
	(x"3cd60000", x"49f30000", x"808e0036", x"aa0a1800", x"89824fd7", x"ec4e516d", x"de1e3a21", x"bbbdaed9", x"68ba0000", x"a0be0000", x"01410031", x"eeea2000", x"bc3a7856", x"a8a5bb57", x"7275e2f2", x"c93a72c5"),
	(x"64950000", x"c98d0000", x"f8bd0037", x"6c612000", x"6eb5130b", x"95e36eb0", x"726dc44e", x"81f9d768", x"75e00000", x"8bcc0000", x"49cc0031", x"418b3800", x"99f15693", x"60dc0487", x"f3d7e6db", x"d74f4463"),
	(x"52500000", x"29540000", x"6a61004e", x"f0ff0000", x"9a317eec", x"452341ce", x"cf568fe5", x"5303130f", x"538d0000", x"a9fc0000", x"9ef70006", x"56ff0000", x"0ae4004e", x"92c5cdf9", x"a9444018", x"7f975691"),
	(x"0a130000", x"a92a0000", x"1252004f", x"36943800", x"7d062230", x"3c8e7e13", x"6325718a", x"69476abe", x"4ed70000", x"828e0000", x"d67a0006", x"f99e1800", x"2f2f2e8b", x"5abc7229", x"28e64431", x"61e26037"),
	(x"4f0a0000", x"02260000", x"22ec004e", x"5f9e1800", x"bffa5029", x"8d5afe1e", x"4ef48bcc", x"4d7625a9", x"16940000", x"02f00000", x"ae490007", x"3ff52000", x"c8187257", x"23114df4", x"8495ba5e", x"5ba61986"),
	(x"17490000", x"82580000", x"5adf004f", x"99f52000", x"58cd0cf5", x"f4f7c1c3", x"e28775a3", x"77325c18", x"0bce0000", x"29820000", x"e6c40007", x"90943800", x"edd35c92", x"eb68f224", x"0537be77", x"45d32f20"),
	(x"f76b0000", x"3d720000", x"24510050", x"8c510000", x"15af7339", x"3dfcebf3", x"3867e73d", x"58185a49", x"54600000", x"1bac0000", x"1983000c", x"c1f20000", x"499623e0", x"da02a35d", x"5d3c223a", x"efe2e75f"),
	(x"af280000", x"bd0c0000", x"5c620051", x"4a3a3800", x"f2982fe5", x"4451d42e", x"94141952", x"625c23f8", x"493a0000", x"30de0000", x"510e000c", x"6e931800", x"6c5d0d25", x"127b1c8d", x"dc9e2613", x"f197d1f9"),
	(x"ea310000", x"16000000", x"6cdc0050", x"23301800", x"30645dfc", x"f5855423", x"b9c5e314", x"466d6cef", x"11790000", x"b0a00000", x"293d000d", x"a8f82000", x"8b6a51f9", x"6bd62350", x"70edd87c", x"cbd3a848"),
	(x"b2720000", x"967e0000", x"14ef0051", x"e55b2000", x"d7530120", x"8c286bfe", x"15b61d7b", x"7c29155e", x"0c230000", x"9bd20000", x"61b0000d", x"07993800", x"aea17f3c", x"a3af9c80", x"f14fdc55", x"d5a69eee"),
	(x"55bd0000", x"9b040000", x"ed150044", x"67f20000", x"d9435d42", x"0de42f6a", x"3b2eedc7", x"c376a2c1", x"f15b0000", x"0f8a0000", x"57b30012", x"bd5c0000", x"c6082e35", x"a2dd0960", x"aa0d4ae2", x"e4f9ae19"),
	(x"0dfe0000", x"1b7a0000", x"95260045", x"a1993800", x"3e74019e", x"744910b7", x"975d13a8", x"f932db70", x"ec010000", x"24f80000", x"1f3e0012", x"123d1800", x"e3c300f0", x"6aa4b6b0", x"2baf4ecb", x"fa8c98bf"),
	(x"48e70000", x"b0760000", x"a5980044", x"c8931800", x"fc887387", x"c59d90ba", x"ba8ce9ee", x"dd039467", x"b4420000", x"a4860000", x"670d0013", x"d4562000", x"04f45c2c", x"1309896d", x"87dcb0a4", x"c0c8e10e"),
	(x"10a40000", x"30080000", x"ddab0045", x"0ef82000", x"1bbf2f5b", x"bc30af67", x"16ff1781", x"e747edd6", x"a9180000", x"8ff40000", x"2f800013", x"7b373800", x"213f72e9", x"db7036bd", x"067eb48d", x"debdd7a8"),
	(x"f0860000", x"8f220000", x"a325005a", x"1b5c0000", x"56dd5097", x"753b8557", x"cc1f851f", x"c86deb87", x"f6b60000", x"bdda0000", x"d0c70018", x"2a510000", x"857a0d9b", x"ea1a67c4", x"5e7528c0", x"748c1fd7"),
	(x"a8c50000", x"0f5c0000", x"db16005b", x"dd373800", x"b1ea0c4b", x"0c96ba8a", x"606c7b70", x"f2299236", x"ebec0000", x"96a80000", x"984a0018", x"85301800", x"a0b1235e", x"2263d814", x"dfd72ce9", x"6af92971"),
	(x"eddc0000", x"a4500000", x"eba8005a", x"b43d1800", x"73167e52", x"bd423a87", x"4dbd8136", x"d618dd21", x"b3af0000", x"16d60000", x"e0790019", x"435b2000", x"47867f82", x"5bcee7c9", x"73a4d286", x"50bd50c0"),
	(x"b59f0000", x"242e0000", x"939b005b", x"72562000", x"9421228e", x"c4ef055a", x"e1ce7f59", x"ec5ca490", x"aef50000", x"3da40000", x"a8f40019", x"ec3a3800", x"624d5147", x"93b75819", x"f206d6af", x"4ec86666"),
	(x"dac80000", x"36c00000", x"15ae0060", x"0bb10000", x"6b697976", x"248dd0a9", x"67c3ff89", x"b513679b", x"584f0000", x"729f0000", x"e07f000a", x"43790000", x"9b1948bd", x"e74476ba", x"5d240486", x"a72142f2"),
	(x"828b0000", x"b6be0000", x"6d9d0061", x"cdda3800", x"8c5e25aa", x"5d20ef74", x"cbb001e6", x"8f571e2a", x"45150000", x"59ed0000", x"a8f2000a", x"ec181800", x"bed26678", x"2f3dc96a", x"dc8600af", x"b9547454"),
	(x"c7920000", x"1db20000", x"5d230060", x"a4d01800", x"4ea257b3", x"ecf46f79", x"e661fba0", x"ab66513d", x"1d560000", x"d9930000", x"d0c1000b", x"2a732000", x"59e53aa4", x"5690f6b7", x"70f5fec0", x"83100de5"),
	(x"9fd10000", x"9dcc0000", x"25100061", x"62bb2000", x"a9950b6f", x"955950a4", x"4a1205cf", x"9122288c", x"000c0000", x"f2e10000", x"984c000b", x"85123800", x"7c2e1461", x"9ee94967", x"f157fae9", x"9d653b43"),
	(x"7ff30000", x"22e60000", x"5b9e007e", x"771f0000", x"e4f774a3", x"5c527a94", x"90f29751", x"be082edd", x"5fa20000", x"c0cf0000", x"670b0000", x"d4740000", x"d86b6b13", x"af83181e", x"a95c66a4", x"3754f33c"),
	(x"27b00000", x"a2980000", x"23ad007f", x"b1743800", x"03c0287f", x"25ff4549", x"3c81693e", x"844c576c", x"42f80000", x"ebbd0000", x"2f860000", x"7b151800", x"fda045d6", x"67faa7ce", x"28fe628d", x"2921c59a"),
	(x"62a90000", x"09940000", x"1313007e", x"d87e1800", x"c13c5a66", x"942bc544", x"11509378", x"a07d187b", x"1abb0000", x"6bc30000", x"57b50001", x"bd7e2000", x"1a97190a", x"1e579813", x"848d9ce2", x"1365bc2b"),
	(x"3aea0000", x"89ea0000", x"6b20007f", x"1e152000", x"260b06ba", x"ed86fa99", x"bd236d17", x"9a3961ca", x"07e10000", x"40b10000", x"1f380001", x"121f3800", x"3f5c37cf", x"d62e27c3", x"052f98cb", x"0d108a8d"),
	(x"dd250000", x"84900000", x"92da006a", x"9cbc0000", x"281b5ad8", x"6c4abe0d", x"93bb9dab", x"2566d655", x"fa990000", x"d4e90000", x"293b001e", x"a8da0000", x"57f566c6", x"d75cb223", x"5e6d0e7c", x"3c4fba7a"),
	(x"85660000", x"04ee0000", x"eae9006b", x"5ad73800", x"cf2c0604", x"15e781d0", x"3fc863c4", x"1f22afe4", x"e7c30000", x"ff9b0000", x"61b6001e", x"07bb1800", x"723e4803", x"1f250df3", x"dfcf0a55", x"223a8cdc"),
	(x"c07f0000", x"afe20000", x"da57006a", x"33dd1800", x"0dd0741d", x"a43301dd", x"12199982", x"3b13e0f3", x"bf800000", x"7fe50000", x"1985001f", x"c1d02000", x"950914df", x"6688322e", x"73bcf43a", x"187ef56d"),
	(x"983c0000", x"2f9c0000", x"a264006b", x"f5b62000", x"eae728c1", x"dd9e3e00", x"be6a67ed", x"01579942", x"a2da0000", x"54970000", x"5108001f", x"6eb13800", x"b0c23a1a", x"aef18dfe", x"f21ef013", x"060bc3cb"),
	(x"781e0000", x"90b60000", x"dcea0074", x"e0120000", x"a785570d", x"14951430", x"648af573", x"2e7d9f13", x"fd740000", x"66b90000", x"ae4f0014", x"3fd70000", x"14874568", x"9f9bdc87", x"aa156c5e", x"ac3a0bb4"),
	(x"205d0000", x"10c80000", x"a4d90075", x"26793800", x"40b20bd1", x"6d382bed", x"c8f90b1c", x"1439e6a2", x"e02e0000", x"4dcb0000", x"e6c20014", x"90b61800", x"314c6bad", x"57e26357", x"2bb76877", x"b24f3d12"),
	(x"65440000", x"bbc40000", x"94670074", x"4f731800", x"824e79c8", x"dcecabe0", x"e528f15a", x"3008a9b5", x"b86d0000", x"cdb50000", x"9ef10015", x"56dd2000", x"d67b3771", x"2e4f5c8a", x"87c49618", x"880b44a3"),
	(x"3d070000", x"3bba0000", x"ec540075", x"89182000", x"65792514", x"a541943d", x"495b0f35", x"0a4cd004", x"a5370000", x"e6c70000", x"d67c0015", x"f9bc3800", x"f3b019b4", x"e636e35a", x"06669231", x"967e7205"),
	(x"59920000", x"f2370000", x"14e90042", x"e5790000", x"0bcc361f", x"30a2fa8d", x"3b36cb7b", x"8bb5076c", x"d0d70000", x"6d0b0000", x"9fb00024", x"b8370000", x"6a414f27", x"86eae7dd", x"f5b174ea", x"41313666"),
	(x"01d10000", x"72490000", x"6cda0043", x"23123800", x"ecfb6ac3", x"490fc550", x"97453514", x"b1f17edd", x"cd8d0000", x"46790000", x"d73d0024", x"17561800", x"4f8a61e2", x"4e93580d", x"741370c3", x"5f4400c0"),
	(x"44c80000", x"d9450000", x"5c640042", x"4a181800", x"2e0718da", x"f8db455d", x"ba94cf52", x"95c031ca", x"95ce0000", x"c6070000", x"af0e0025", x"d13d2000", x"a8bd3d3e", x"373e67d0", x"d8608eac", x"65007971"),
	(x"1c8b0000", x"593b0000", x"24570043", x"8c732000", x"c9304406", x"81767a80", x"16e7313d", x"af84487b", x"88940000", x"ed750000", x"e7830025", x"7e5c3800", x"8d7613fb", x"ff47d800", x"59c28a85", x"7b754fd7"),
	(x"fca90000", x"e6110000", x"5ad9005c", x"99d70000", x"84523bca", x"487d50b0", x"cc07a3a3", x"80ae4e2a", x"d73a0000", x"df5b0000", x"18c4002e", x"2f3a0000", x"29336c89", x"ce2d8979", x"01c916c8", x"d14487a8"),
	(x"a4ea0000", x"666f0000", x"22ea005d", x"5fbc3800", x"63656716", x"31d06f6d", x"60745dcc", x"baea379b", x"ca600000", x"f4290000", x"5049002e", x"805b1800", x"0cf8424c", x"065436a9", x"806b12e1", x"cf31b10e"),
	(x"e1f30000", x"cd630000", x"1254005c", x"36b61800", x"a199150f", x"8004ef60", x"4da5a78a", x"9edb788c", x"92230000", x"74570000", x"287a002f", x"46302000", x"ebcf1e90", x"7ff90974", x"2c18ec8e", x"f575c8bf"),
	(x"b9b00000", x"4d1d0000", x"6a67005d", x"f0dd2000", x"46ae49d3", x"f9a9d0bd", x"e1d659e5", x"a49f013d", x"8f790000", x"5f250000", x"60f7002f", x"e9513800", x"ce043055", x"b780b6a4", x"adbae8a7", x"eb00fe19"),
	(x"5e7f0000", x"40670000", x"939d0048", x"72740000", x"48be15b1", x"78659429", x"cf4ea959", x"1bc0b6a2", x"72010000", x"cb7d0000", x"56f40030", x"53940000", x"a6ad615c", x"b6f22344", x"f6f87e10", x"da5fceee"),
	(x"063c0000", x"c0190000", x"ebae0049", x"b41f3800", x"af89496d", x"01c8abf4", x"633d5736", x"2184cf13", x"6f5b0000", x"e00f0000", x"1e790030", x"fcf51800", x"83664f99", x"7e8b9c94", x"775a7a39", x"c42af848"),
	(x"43250000", x"6b150000", x"db100048", x"dd151800", x"6d753b74", x"b01c2bf9", x"4eecad70", x"05b58004", x"37180000", x"60710000", x"664a0031", x"3a9e2000", x"64511345", x"0726a349", x"db298456", x"fe6e81f9"),
	(x"1b660000", x"eb6b0000", x"a3230049", x"1b7e2000", x"8a4267a8", x"c9b11424", x"e29f531f", x"3ff1f9b5", x"2a420000", x"4b030000", x"2ec70031", x"95ff3800", x"419a3d80", x"cf5f1c99", x"5a8b807f", x"e01bb75f"),
	(x"fb440000", x"54410000", x"ddad0056", x"0eda0000", x"c7201864", x"00ba3e14", x"387fc181", x"10dbffe4", x"75ec0000", x"792d0000", x"d180003a", x"c4990000", x"e5df42f2", x"fe354de0", x"02801c32", x"4a2a7f20"),
	(x"a3070000", x"d43f0000", x"a59e0057", x"c8b13800", x"201744b8", x"791701c9", x"940c3fee", x"2a9f8655", x"68b60000", x"525f0000", x"990d003a", x"6bf81800", x"c0146c37", x"364cf230", x"8322181b", x"545f4986"),
	(x"e61e0000", x"7f330000", x"95200056", x"a1bb1800", x"e2eb36a1", x"c8c381c4", x"b9ddc5a8", x"0eaec942", x"30f50000", x"d2210000", x"e13e003b", x"ad932000", x"272330eb", x"4fe1cded", x"2f51e674", x"6e1b3037"),
	(x"be5d0000", x"ff4d0000", x"ed130057", x"67d02000", x"05dc6a7d", x"b16ebe19", x"15ae3bc7", x"34eab0f3", x"2daf0000", x"f9530000", x"a9b3003b", x"02f23800", x"02e81e2e", x"8798723d", x"aef3e25d", x"706e0691"),
	(x"d10a0000", x"eda30000", x"6b26006c", x"1e370000", x"fa943185", x"510c6bea", x"93a3bb17", x"6da573f8", x"db150000", x"b6680000", x"e1380028", x"adb10000", x"fbbc07d4", x"f36b5c9e", x"01d13074", x"99872205"),
	(x"89490000", x"6ddd0000", x"1315006d", x"d85c3800", x"1da36d59", x"28a15437", x"3fd04578", x"57e10a49", x"c64f0000", x"9d1a0000", x"a9b50028", x"02d01800", x"de772911", x"3b12e34e", x"8073345d", x"87f214a3"),
	(x"cc500000", x"c6d10000", x"23ab006c", x"b1561800", x"df5f1f40", x"9975d43a", x"1201bf3e", x"73d0455e", x"9e0c0000", x"1d640000", x"d1860029", x"c4bb2000", x"394075cd", x"42bfdc93", x"2c00ca32", x"bdb66d12"),
	(x"94130000", x"46af0000", x"5b98006d", x"773d2000", x"3868439c", x"e0d8ebe7", x"be724151", x"49943cef", x"83560000", x"36160000", x"990b0029", x"6bda3800", x"1c8b5b08", x"8ac66343", x"ada2ce1b", x"a3c35bb4"),
	(x"74310000", x"f9850000", x"25160072", x"62990000", x"750a3c50", x"29d3c1d7", x"6492d3cf", x"66be3abe", x"dcf80000", x"04380000", x"664c0022", x"3abc0000", x"b8ce247a", x"bbac323a", x"f5a95256", x"09f293cb"),
	(x"2c720000", x"79fb0000", x"5d250073", x"a4f23800", x"923d608c", x"507efe0a", x"c8e12da0", x"5cfa430f", x"c1a20000", x"2f4a0000", x"2ec10022", x"95dd1800", x"9d050abf", x"73d58dea", x"740b567f", x"1787a56d"),
	(x"696b0000", x"d2f70000", x"6d9b0072", x"cdf81800", x"50c11295", x"e1aa7e07", x"e530d7e6", x"78cb0c18", x"99e10000", x"af340000", x"56f20023", x"53b62000", x"7a325663", x"0a78b237", x"d878a810", x"2dc3dcdc"),
	(x"31280000", x"52890000", x"15a80073", x"0b932000", x"b7f64e49", x"980741da", x"49432989", x"428f75a9", x"84bb0000", x"84460000", x"1e7f0023", x"fcd73800", x"5ff978a6", x"c2010de7", x"59daac39", x"33b6ea7a"),
	(x"d6e70000", x"5ff30000", x"ec520066", x"893a0000", x"b9e6122b", x"19cb054e", x"67dbd935", x"fdd0c236", x"79c30000", x"101e0000", x"287c003c", x"46120000", x"375029af", x"c3739807", x"02983a8e", x"02e9da8d"),
	(x"8ea40000", x"df8d0000", x"94610067", x"4f513800", x"5ed14ef7", x"60663a93", x"cba8275a", x"c794bb87", x"64990000", x"3b6c0000", x"60f1003c", x"e9731800", x"129b076a", x"0b0a27d7", x"833a3ea7", x"1c9cec2b"),
	(x"cbbd0000", x"74810000", x"a4df0066", x"265b1800", x"9c2d3cee", x"d1b2ba9e", x"e679dd1c", x"e3a5f490", x"3cda0000", x"bb120000", x"18c2003d", x"2f182000", x"f5ac5bb6", x"72a7180a", x"2f49c0c8", x"26d8959a"),
	(x"93fe0000", x"f4ff0000", x"dcec0067", x"e0302000", x"7b1a6032", x"a81f8543", x"4a0a2373", x"d9e18d21", x"21800000", x"90600000", x"504f003d", x"80793800", x"d0677573", x"badea7da", x"aeebc4e1", x"38ada33c"),
	(x"73dc0000", x"4bd50000", x"a2620078", x"f5940000", x"36781ffe", x"6114af73", x"90eab1ed", x"f6cb8b70", x"7e2e0000", x"a24e0000", x"af080036", x"d11f0000", x"74220a01", x"8bb4f6a3", x"f6e058ac", x"929c6b43"),
	(x"2b9f0000", x"cbab0000", x"da510079", x"33ff3800", x"d14f4322", x"18b990ae", x"3c994f82", x"cc8ff2c1", x"63740000", x"893c0000", x"e7850036", x"7e7e1800", x"51e924c4", x"43cd4973", x"77425c85", x"8ce95de5"),
	(x"6e860000", x"60a70000", x"eaef0078", x"5af51800", x"13b3313b", x"a96d10a3", x"1148b5c4", x"e8bebdd6", x"3b370000", x"09420000", x"9fb60037", x"b8152000", x"b6de7818", x"3a6076ae", x"db31a2ea", x"b6ad2454"),
	(x"36c50000", x"e0d90000", x"92dc0079", x"9c9e2000", x"f4846de7", x"d0c02f7e", x"bd3b4bab", x"d2fac467", x"266d0000", x"22300000", x"d73b0037", x"17743800", x"931556dd", x"f219c97e", x"5a93a6c3", x"a8d812f2"),
	(x"538d0000", x"a9fc0000", x"9ef70006", x"56ff0000", x"0ae4004e", x"92c5cdf9", x"a9444018", x"7f975691", x"01dd0000", x"80a80000", x"f4960048", x"a6000000", x"90d57ea2", x"d7e68c37", x"6612cffd", x"2c94459e"),
	(x"0bce0000", x"29820000", x"e6c40007", x"90943800", x"edd35c92", x"eb68f224", x"0537be77", x"45d32f20", x"1c870000", x"abda0000", x"bc1b0048", x"09611800", x"b51e5067", x"1f9f33e7", x"e7b0cbd4", x"32e17338"),
	(x"4ed70000", x"828e0000", x"d67a0006", x"f99e1800", x"2f2f2e8b", x"5abc7229", x"28e64431", x"61e26037", x"44c40000", x"2ba40000", x"c4280049", x"cf0a2000", x"52290cbb", x"66320c3a", x"4bc335bb", x"08a50a89"),
	(x"16940000", x"02f00000", x"ae490007", x"3ff52000", x"c8187257", x"23114df4", x"8495ba5e", x"5ba61986", x"599e0000", x"00d60000", x"8ca50049", x"606b3800", x"77e2227e", x"ae4bb3ea", x"ca613192", x"16d03c2f"),
	(x"f6b60000", x"bdda0000", x"d0c70018", x"2a510000", x"857a0d9b", x"ea1a67c4", x"5e7528c0", x"748c1fd7", x"06300000", x"32f80000", x"73e20042", x"310d0000", x"d3a75d0c", x"9f21e293", x"926aaddf", x"bce1f450"),
	(x"aef50000", x"3da40000", x"a8f40019", x"ec3a3800", x"624d5147", x"93b75819", x"f206d6af", x"4ec86666", x"1b6a0000", x"198a0000", x"3b6f0042", x"9e6c1800", x"f66c73c9", x"57585d43", x"13c8a9f6", x"a294c2f6"),
	(x"ebec0000", x"96a80000", x"984a0018", x"85301800", x"a0b1235e", x"2263d814", x"dfd72ce9", x"6af92971", x"43290000", x"99f40000", x"435c0043", x"58072000", x"115b2f15", x"2ef5629e", x"bfbb5799", x"98d0bb47"),
	(x"b3af0000", x"16d60000", x"e0790019", x"435b2000", x"47867f82", x"5bcee7c9", x"73a4d286", x"50bd50c0", x"5e730000", x"b2860000", x"0bd10043", x"f7663800", x"349001d0", x"e68cdd4e", x"3e1953b0", x"86a58de1"),
	(x"54600000", x"1bac0000", x"1983000c", x"c1f20000", x"499623e0", x"da02a35d", x"5d3c223a", x"efe2e75f", x"a30b0000", x"26de0000", x"3dd2005c", x"4da30000", x"5c3950d9", x"e7fe48ae", x"655bc507", x"b7fabd16"),
	(x"0c230000", x"9bd20000", x"61b0000d", x"07993800", x"aea17f3c", x"a3af9c80", x"f14fdc55", x"d5a69eee", x"be510000", x"0dac0000", x"755f005c", x"e2c21800", x"79f27e1c", x"2f87f77e", x"e4f9c12e", x"a98f8bb0"),
	(x"493a0000", x"30de0000", x"510e000c", x"6e931800", x"6c5d0d25", x"127b1c8d", x"dc9e2613", x"f197d1f9", x"e6120000", x"8dd20000", x"0d6c005d", x"24a92000", x"9ec522c0", x"562ac8a3", x"488a3f41", x"93cbf201"),
	(x"11790000", x"b0a00000", x"293d000d", x"a8f82000", x"8b6a51f9", x"6bd62350", x"70edd87c", x"cbd3a848", x"fb480000", x"a6a00000", x"45e1005d", x"8bc83800", x"bb0e0c05", x"9e537773", x"c9283b68", x"8dbec4a7"),
	(x"f15b0000", x"0f8a0000", x"57b30012", x"bd5c0000", x"c6082e35", x"a2dd0960", x"aa0d4ae2", x"e4f9ae19", x"a4e60000", x"948e0000", x"baa60056", x"daae0000", x"1f4b7377", x"af39260a", x"9123a725", x"278f0cd8"),
	(x"a9180000", x"8ff40000", x"2f800013", x"7b373800", x"213f72e9", x"db7036bd", x"067eb48d", x"debdd7a8", x"b9bc0000", x"bffc0000", x"f22b0056", x"75cf1800", x"3a805db2", x"674099da", x"1081a30c", x"39fa3a7e"),
	(x"ec010000", x"24f80000", x"1f3e0012", x"123d1800", x"e3c300f0", x"6aa4b6b0", x"2baf4ecb", x"fa8c98bf", x"e1ff0000", x"3f820000", x"8a180057", x"b3a42000", x"ddb7016e", x"1eeda607", x"bcf25d63", x"03be43cf"),
	(x"b4420000", x"a4860000", x"670d0013", x"d4562000", x"04f45c2c", x"1309896d", x"87dcb0a4", x"c0c8e10e", x"fca50000", x"14f00000", x"c2950057", x"1cc53800", x"f87c2fab", x"d69419d7", x"3d50594a", x"1dcb7569"),
	(x"db150000", x"b6680000", x"e1380028", x"adb10000", x"fbbc07d4", x"f36b5c9e", x"01d13074", x"99872205", x"0a1f0000", x"5bcb0000", x"8a1e0044", x"b3860000", x"01283651", x"a2673774", x"92728b63", x"f42251fd"),
	(x"83560000", x"36160000", x"990b0029", x"6bda3800", x"1c8b5b08", x"8ac66343", x"ada2ce1b", x"a3c35bb4", x"17450000", x"70b90000", x"c2930044", x"1ce71800", x"24e31894", x"6a1e88a4", x"13d08f4a", x"ea57675b"),
	(x"c64f0000", x"9d1a0000", x"a9b50028", x"02d01800", x"de772911", x"3b12e34e", x"8073345d", x"87f214a3", x"4f060000", x"f0c70000", x"baa00045", x"da8c2000", x"c3d44448", x"13b3b779", x"bfa37125", x"d0131eea"),
	(x"9e0c0000", x"1d640000", x"d1860029", x"c4bb2000", x"394075cd", x"42bfdc93", x"2c00ca32", x"bdb66d12", x"525c0000", x"dbb50000", x"f22d0045", x"75ed3800", x"e61f6a8d", x"dbca08a9", x"3e01750c", x"ce66284c"),
	(x"7e2e0000", x"a24e0000", x"af080036", x"d11f0000", x"74220a01", x"8bb4f6a3", x"f6e058ac", x"929c6b43", x"0df20000", x"e99b0000", x"0d6a004e", x"248b0000", x"425a15ff", x"eaa059d0", x"660ae941", x"6457e033"),
	(x"266d0000", x"22300000", x"d73b0037", x"17743800", x"931556dd", x"f219c97e", x"5a93a6c3", x"a8d812f2", x"10a80000", x"c2e90000", x"45e7004e", x"8bea1800", x"67913b3a", x"22d9e600", x"e7a8ed68", x"7a22d695"),
	(x"63740000", x"893c0000", x"e7850036", x"7e7e1800", x"51e924c4", x"43cd4973", x"77425c85", x"8ce95de5", x"48eb0000", x"42970000", x"3dd4004f", x"4d812000", x"80a667e6", x"5b74d9dd", x"4bdb1307", x"4066af24"),
	(x"3b370000", x"09420000", x"9fb60037", x"b8152000", x"b6de7818", x"3a6076ae", x"db31a2ea", x"b6ad2454", x"55b10000", x"69e50000", x"7559004f", x"e2e03800", x"a56d4923", x"930d660d", x"ca79172e", x"5e139982"),
	(x"dcf80000", x"04380000", x"664c0022", x"3abc0000", x"b8ce247a", x"bbac323a", x"f5a95256", x"09f293cb", x"a8c90000", x"fdbd0000", x"435a0050", x"58250000", x"cdc4182a", x"927ff3ed", x"913b8199", x"6f4ca975"),
	(x"84bb0000", x"84460000", x"1e7f0023", x"fcd73800", x"5ff978a6", x"c2010de7", x"59daac39", x"33b6ea7a", x"b5930000", x"d6cf0000", x"0bd70050", x"f7441800", x"e80f36ef", x"5a064c3d", x"109985b0", x"71399fd3"),
	(x"c1a20000", x"2f4a0000", x"2ec10022", x"95dd1800", x"9d050abf", x"73d58dea", x"740b567f", x"1787a56d", x"edd00000", x"56b10000", x"73e40051", x"312f2000", x"0f386a33", x"23ab73e0", x"bcea7bdf", x"4b7de662"),
	(x"99e10000", x"af340000", x"56f20023", x"53b62000", x"7a325663", x"0a78b237", x"d878a810", x"2dc3dcdc", x"f08a0000", x"7dc30000", x"3b690051", x"9e4e3800", x"2af344f6", x"ebd2cc30", x"3d487ff6", x"5508d0c4"),
	(x"79c30000", x"101e0000", x"287c003c", x"46120000", x"375029af", x"c3739807", x"02983a8e", x"02e9da8d", x"af240000", x"4fed0000", x"c42e005a", x"cf280000", x"8eb63b84", x"dab89d49", x"6543e3bb", x"ff3918bb"),
	(x"21800000", x"90600000", x"504f003d", x"80793800", x"d0677573", x"badea7da", x"aeebc4e1", x"38ada33c", x"b27e0000", x"649f0000", x"8ca3005a", x"60491800", x"ab7d1541", x"12c12299", x"e4e1e792", x"e14c2e1d"),
	(x"64990000", x"3b6c0000", x"60f1003c", x"e9731800", x"129b076a", x"0b0a27d7", x"833a3ea7", x"1c9cec2b", x"ea3d0000", x"e4e10000", x"f490005b", x"a6222000", x"4c4a499d", x"6b6c1d44", x"489219fd", x"db0857ac"),
	(x"3cda0000", x"bb120000", x"18c2003d", x"2f182000", x"f5ac5bb6", x"72a7180a", x"2f49c0c8", x"26d8959a", x"f7670000", x"cf930000", x"bc1d005b", x"09433800", x"69816758", x"a315a294", x"c9301dd4", x"c57d610a"),
	(x"584f0000", x"729f0000", x"e07f000a", x"43790000", x"9b1948bd", x"e74476ba", x"5d240486", x"a72142f2", x"82870000", x"445f0000", x"f5d1006a", x"48c80000", x"f07031cb", x"c3c9a613", x"3ae7fb0f", x"12322569"),
	(x"000c0000", x"f2e10000", x"984c000b", x"85123800", x"7c2e1461", x"9ee94967", x"f157fae9", x"9d653b43", x"9fdd0000", x"6f2d0000", x"bd5c006a", x"e7a91800", x"d5bb1f0e", x"0bb019c3", x"bb45ff26", x"0c4713cf"),
	(x"45150000", x"59ed0000", x"a8f2000a", x"ec181800", x"bed26678", x"2f3dc96a", x"dc8600af", x"b9547454", x"c79e0000", x"ef530000", x"c56f006b", x"21c22000", x"328c43d2", x"721d261e", x"17360149", x"36036a7e"),
	(x"1d560000", x"d9930000", x"d0c1000b", x"2a732000", x"59e53aa4", x"5690f6b7", x"70f5fec0", x"83100de5", x"dac40000", x"c4210000", x"8de2006b", x"8ea33800", x"17476d17", x"ba6499ce", x"96940560", x"28765cd8"),
	(x"fd740000", x"66b90000", x"ae4f0014", x"3fd70000", x"14874568", x"9f9bdc87", x"aa156c5e", x"ac3a0bb4", x"856a0000", x"f60f0000", x"72a50060", x"dfc50000", x"b3021265", x"8b0ec8b7", x"ce9f992d", x"824794a7"),
	(x"a5370000", x"e6c70000", x"d67c0015", x"f9bc3800", x"f3b019b4", x"e636e35a", x"06669231", x"967e7205", x"98300000", x"dd7d0000", x"3a280060", x"70a41800", x"96c93ca0", x"43777767", x"4f3d9d04", x"9c32a201"),
	(x"e02e0000", x"4dcb0000", x"e6c20014", x"90b61800", x"314c6bad", x"57e26357", x"2bb76877", x"b24f3d12", x"c0730000", x"5d030000", x"421b0061", x"b6cf2000", x"71fe607c", x"3ada48ba", x"e34e636b", x"a676dbb0"),
	(x"b86d0000", x"cdb50000", x"9ef10015", x"56dd2000", x"d67b3771", x"2e4f5c8a", x"87c49618", x"880b44a3", x"dd290000", x"76710000", x"0a960061", x"19ae3800", x"54354eb9", x"f2a3f76a", x"62ec6742", x"b803ed16"),
	(x"5fa20000", x"c0cf0000", x"670b0000", x"d4740000", x"d86b6b13", x"af83181e", x"a95c66a4", x"3754f33c", x"20510000", x"e2290000", x"3c95007e", x"a36b0000", x"3c9c1fb0", x"f3d1628a", x"39aef1f5", x"895cdde1"),
	(x"07e10000", x"40b10000", x"1f380001", x"121f3800", x"3f5c37cf", x"d62e27c3", x"052f98cb", x"0d108a8d", x"3d0b0000", x"c95b0000", x"7418007e", x"0c0a1800", x"19573175", x"3ba8dd5a", x"b80cf5dc", x"9729eb47"),
	(x"42f80000", x"ebbd0000", x"2f860000", x"7b151800", x"fda045d6", x"67faa7ce", x"28fe628d", x"2921c59a", x"65480000", x"49250000", x"0c2b007f", x"ca612000", x"fe606da9", x"4205e287", x"147f0bb3", x"ad6d92f6"),
	(x"1abb0000", x"6bc30000", x"57b50001", x"bd7e2000", x"1a97190a", x"1e579813", x"848d9ce2", x"1365bc2b", x"78120000", x"62570000", x"44a6007f", x"65003800", x"dbab436c", x"8a7c5d57", x"95dd0f9a", x"b318a450"),
	(x"fa990000", x"d4e90000", x"293b001e", x"a8da0000", x"57f566c6", x"d75cb223", x"5e6d0e7c", x"3c4fba7a", x"27bc0000", x"50790000", x"bbe10074", x"34660000", x"7fee3c1e", x"bb160c2e", x"cdd693d7", x"19296c2f"),
	(x"a2da0000", x"54970000", x"5108001f", x"6eb13800", x"b0c23a1a", x"aef18dfe", x"f21ef013", x"060bc3cb", x"3ae60000", x"7b0b0000", x"f36c0074", x"9b071800", x"5a2512db", x"736fb3fe", x"4c7497fe", x"075c5a89"),
	(x"e7c30000", x"ff9b0000", x"61b6001e", x"07bb1800", x"723e4803", x"1f250df3", x"dfcf0a55", x"223a8cdc", x"62a50000", x"fb750000", x"8b5f0075", x"5d6c2000", x"bd124e07", x"0ac28c23", x"e0076991", x"3d182338"),
	(x"bf800000", x"7fe50000", x"1985001f", x"c1d02000", x"950914df", x"6688322e", x"73bcf43a", x"187ef56d", x"7fff0000", x"d0070000", x"c3d20075", x"f20d3800", x"98d960c2", x"c2bb33f3", x"61a56db8", x"236d159e"),
	(x"d0d70000", x"6d0b0000", x"9fb00024", x"b8370000", x"6a414f27", x"86eae7dd", x"f5b174ea", x"41313666", x"89450000", x"9f3c0000", x"8b590066", x"5d4e0000", x"618d7938", x"b6481d50", x"ce87bf91", x"ca84310a"),
	(x"88940000", x"ed750000", x"e7830025", x"7e5c3800", x"8d7613fb", x"ff47d800", x"59c28a85", x"7b754fd7", x"941f0000", x"b44e0000", x"c3d40066", x"f22f1800", x"444657fd", x"7e31a280", x"4f25bbb8", x"d4f107ac"),
	(x"cd8d0000", x"46790000", x"d73d0024", x"17561800", x"4f8a61e2", x"4e93580d", x"741370c3", x"5f4400c0", x"cc5c0000", x"34300000", x"bbe70067", x"34442000", x"a3710b21", x"079c9d5d", x"e35645d7", x"eeb57e1d"),
	(x"95ce0000", x"c6070000", x"af0e0025", x"d13d2000", x"a8bd3d3e", x"373e67d0", x"d8608eac", x"65007971", x"d1060000", x"1f420000", x"f36a0067", x"9b253800", x"86ba25e4", x"cfe5228d", x"62f441fe", x"f0c048bb"),
	(x"75ec0000", x"792d0000", x"d180003a", x"c4990000", x"e5df42f2", x"fe354de0", x"02801c32", x"4a2a7f20", x"8ea80000", x"2d6c0000", x"0c2d006c", x"ca430000", x"22ff5a96", x"fe8f73f4", x"3affddb3", x"5af180c4"),
	(x"2daf0000", x"f9530000", x"a9b3003b", x"02f23800", x"02e81e2e", x"8798723d", x"aef3e25d", x"706e0691", x"93f20000", x"061e0000", x"44a0006c", x"65221800", x"07347453", x"36f6cc24", x"bb5dd99a", x"4484b662"),
	(x"68b60000", x"525f0000", x"990d003a", x"6bf81800", x"c0146c37", x"364cf230", x"8322181b", x"545f4986", x"cbb10000", x"86600000", x"3c93006d", x"a3492000", x"e003288f", x"4f5bf3f9", x"172e27f5", x"7ec0cfd3"),
	(x"30f50000", x"d2210000", x"e13e003b", x"ad932000", x"272330eb", x"4fe1cded", x"2f51e674", x"6e1b3037", x"d6eb0000", x"ad120000", x"741e006d", x"0c283800", x"c5c8064a", x"87224c29", x"968c23dc", x"60b5f975"),
	(x"d73a0000", x"df5b0000", x"18c4002e", x"2f3a0000", x"29336c89", x"ce2d8979", x"01c916c8", x"d14487a8", x"2b930000", x"394a0000", x"421d0072", x"b6ed0000", x"ad615743", x"8650d9c9", x"cdceb56b", x"51eac982"),
	(x"8f790000", x"5f250000", x"60f7002f", x"e9513800", x"ce043055", x"b780b6a4", x"adbae8a7", x"eb00fe19", x"36c90000", x"12380000", x"0a900072", x"198c1800", x"88aa7986", x"4e296619", x"4c6cb142", x"4f9fff24"),
	(x"ca600000", x"f4290000", x"5049002e", x"805b1800", x"0cf8424c", x"065436a9", x"806b12e1", x"cf31b10e", x"6e8a0000", x"92460000", x"72a30073", x"dfe72000", x"6f9d255a", x"378459c4", x"e01f4f2d", x"75db8695"),
	(x"92230000", x"74570000", x"287a002f", x"46302000", x"ebcf1e90", x"7ff90974", x"2c18ec8e", x"f575c8bf", x"73d00000", x"b9340000", x"3a2e0073", x"70863800", x"4a560b9f", x"fffde614", x"61bd4b04", x"6baeb033"),
	(x"72010000", x"cb7d0000", x"56f40030", x"53940000", x"a6ad615c", x"b6f22344", x"f6f87e10", x"da5fceee", x"2c7e0000", x"8b1a0000", x"c5690078", x"21e00000", x"ee1374ed", x"ce97b76d", x"39b6d749", x"c19f784c"),
	(x"2a420000", x"4b030000", x"2ec70031", x"95ff3800", x"419a3d80", x"cf5f1c99", x"5a8b807f", x"e01bb75f", x"31240000", x"a0680000", x"8de40078", x"8e811800", x"cbd85a28", x"06ee08bd", x"b814d360", x"dfea4eea"),
	(x"6f5b0000", x"e00f0000", x"1e790030", x"fcf51800", x"83664f99", x"7e8b9c94", x"775a7a39", x"c42af848", x"69670000", x"20160000", x"f5d70079", x"48ea2000", x"2cef06f4", x"7f433760", x"14672d0f", x"e5ae375b"),
	(x"37180000", x"60710000", x"664a0031", x"3a9e2000", x"64511345", x"0726a349", x"db298456", x"fe6e81f9", x"743d0000", x"0b640000", x"bd5a0079", x"e78b3800", x"09242831", x"b73a88b0", x"95c52926", x"fbdb01fd"),
	(x"01dd0000", x"80a80000", x"f4960048", x"a6000000", x"90d57ea2", x"d7e68c37", x"6612cffd", x"2c94459e", x"52500000", x"29540000", x"6a61004e", x"f0ff0000", x"9a317eec", x"452341ce", x"cf568fe5", x"5303130f"),
	(x"599e0000", x"00d60000", x"8ca50049", x"606b3800", x"77e2227e", x"ae4bb3ea", x"ca613192", x"16d03c2f", x"4f0a0000", x"02260000", x"22ec004e", x"5f9e1800", x"bffa5029", x"8d5afe1e", x"4ef48bcc", x"4d7625a9"),
	(x"1c870000", x"abda0000", x"bc1b0048", x"09611800", x"b51e5067", x"1f9f33e7", x"e7b0cbd4", x"32e17338", x"17490000", x"82580000", x"5adf004f", x"99f52000", x"58cd0cf5", x"f4f7c1c3", x"e28775a3", x"77325c18"),
	(x"44c40000", x"2ba40000", x"c4280049", x"cf0a2000", x"52290cbb", x"66320c3a", x"4bc335bb", x"08a50a89", x"0a130000", x"a92a0000", x"1252004f", x"36943800", x"7d062230", x"3c8e7e13", x"6325718a", x"69476abe"),
	(x"a4e60000", x"948e0000", x"baa60056", x"daae0000", x"1f4b7377", x"af39260a", x"9123a725", x"278f0cd8", x"55bd0000", x"9b040000", x"ed150044", x"67f20000", x"d9435d42", x"0de42f6a", x"3b2eedc7", x"c376a2c1"),
	(x"fca50000", x"14f00000", x"c2950057", x"1cc53800", x"f87c2fab", x"d69419d7", x"3d50594a", x"1dcb7569", x"48e70000", x"b0760000", x"a5980044", x"c8931800", x"fc887387", x"c59d90ba", x"ba8ce9ee", x"dd039467"),
	(x"b9bc0000", x"bffc0000", x"f22b0056", x"75cf1800", x"3a805db2", x"674099da", x"1081a30c", x"39fa3a7e", x"10a40000", x"30080000", x"ddab0045", x"0ef82000", x"1bbf2f5b", x"bc30af67", x"16ff1781", x"e747edd6"),
	(x"e1ff0000", x"3f820000", x"8a180057", x"b3a42000", x"ddb7016e", x"1eeda607", x"bcf25d63", x"03be43cf", x"0dfe0000", x"1b7a0000", x"95260045", x"a1993800", x"3e74019e", x"744910b7", x"975d13a8", x"f932db70"),
	(x"06300000", x"32f80000", x"73e20042", x"310d0000", x"d3a75d0c", x"9f21e293", x"926aaddf", x"bce1f450", x"f0860000", x"8f220000", x"a325005a", x"1b5c0000", x"56dd5097", x"753b8557", x"cc1f851f", x"c86deb87"),
	(x"5e730000", x"b2860000", x"0bd10043", x"f7663800", x"349001d0", x"e68cdd4e", x"3e1953b0", x"86a58de1", x"eddc0000", x"a4500000", x"eba8005a", x"b43d1800", x"73167e52", x"bd423a87", x"4dbd8136", x"d618dd21"),
	(x"1b6a0000", x"198a0000", x"3b6f0042", x"9e6c1800", x"f66c73c9", x"57585d43", x"13c8a9f6", x"a294c2f6", x"b59f0000", x"242e0000", x"939b005b", x"72562000", x"9421228e", x"c4ef055a", x"e1ce7f59", x"ec5ca490"),
	(x"43290000", x"99f40000", x"435c0043", x"58072000", x"115b2f15", x"2ef5629e", x"bfbb5799", x"98d0bb47", x"a8c50000", x"0f5c0000", x"db16005b", x"dd373800", x"b1ea0c4b", x"0c96ba8a", x"606c7b70", x"f2299236"),
	(x"a30b0000", x"26de0000", x"3dd2005c", x"4da30000", x"5c3950d9", x"e7fe48ae", x"655bc507", x"b7fabd16", x"f76b0000", x"3d720000", x"24510050", x"8c510000", x"15af7339", x"3dfcebf3", x"3867e73d", x"58185a49"),
	(x"fb480000", x"a6a00000", x"45e1005d", x"8bc83800", x"bb0e0c05", x"9e537773", x"c9283b68", x"8dbec4a7", x"ea310000", x"16000000", x"6cdc0050", x"23301800", x"30645dfc", x"f5855423", x"b9c5e314", x"466d6cef"),
	(x"be510000", x"0dac0000", x"755f005c", x"e2c21800", x"79f27e1c", x"2f87f77e", x"e4f9c12e", x"a98f8bb0", x"b2720000", x"967e0000", x"14ef0051", x"e55b2000", x"d7530120", x"8c286bfe", x"15b61d7b", x"7c29155e"),
	(x"e6120000", x"8dd20000", x"0d6c005d", x"24a92000", x"9ec522c0", x"562ac8a3", x"488a3f41", x"93cbf201", x"af280000", x"bd0c0000", x"5c620051", x"4a3a3800", x"f2982fe5", x"4451d42e", x"94141952", x"625c23f8"),
	(x"89450000", x"9f3c0000", x"8b590066", x"5d4e0000", x"618d7938", x"b6481d50", x"ce87bf91", x"ca84310a", x"59920000", x"f2370000", x"14e90042", x"e5790000", x"0bcc361f", x"30a2fa8d", x"3b36cb7b", x"8bb5076c"),
	(x"d1060000", x"1f420000", x"f36a0067", x"9b253800", x"86ba25e4", x"cfe5228d", x"62f441fe", x"f0c048bb", x"44c80000", x"d9450000", x"5c640042", x"4a181800", x"2e0718da", x"f8db455d", x"ba94cf52", x"95c031ca"),
	(x"941f0000", x"b44e0000", x"c3d40066", x"f22f1800", x"444657fd", x"7e31a280", x"4f25bbb8", x"d4f107ac", x"1c8b0000", x"593b0000", x"24570043", x"8c732000", x"c9304406", x"81767a80", x"16e7313d", x"af84487b"),
	(x"cc5c0000", x"34300000", x"bbe70067", x"34442000", x"a3710b21", x"079c9d5d", x"e35645d7", x"eeb57e1d", x"01d10000", x"72490000", x"6cda0043", x"23123800", x"ecfb6ac3", x"490fc550", x"97453514", x"b1f17edd"),
	(x"2c7e0000", x"8b1a0000", x"c5690078", x"21e00000", x"ee1374ed", x"ce97b76d", x"39b6d749", x"c19f784c", x"5e7f0000", x"40670000", x"939d0048", x"72740000", x"48be15b1", x"78659429", x"cf4ea959", x"1bc0b6a2"),
	(x"743d0000", x"0b640000", x"bd5a0079", x"e78b3800", x"09242831", x"b73a88b0", x"95c52926", x"fbdb01fd", x"43250000", x"6b150000", x"db100048", x"dd151800", x"6d753b74", x"b01c2bf9", x"4eecad70", x"05b58004"),
	(x"31240000", x"a0680000", x"8de40078", x"8e811800", x"cbd85a28", x"06ee08bd", x"b814d360", x"dfea4eea", x"1b660000", x"eb6b0000", x"a3230049", x"1b7e2000", x"8a4267a8", x"c9b11424", x"e29f531f", x"3ff1f9b5"),
	(x"69670000", x"20160000", x"f5d70079", x"48ea2000", x"2cef06f4", x"7f433760", x"14672d0f", x"e5ae375b", x"063c0000", x"c0190000", x"ebae0049", x"b41f3800", x"af89496d", x"01c8abf4", x"633d5736", x"2184cf13"),
	(x"8ea80000", x"2d6c0000", x"0c2d006c", x"ca430000", x"22ff5a96", x"fe8f73f4", x"3affddb3", x"5af180c4", x"fb440000", x"54410000", x"ddad0056", x"0eda0000", x"c7201864", x"00ba3e14", x"387fc181", x"10dbffe4"),
	(x"d6eb0000", x"ad120000", x"741e006d", x"0c283800", x"c5c8064a", x"87224c29", x"968c23dc", x"60b5f975", x"e61e0000", x"7f330000", x"95200056", x"a1bb1800", x"e2eb36a1", x"c8c381c4", x"b9ddc5a8", x"0eaec942"),
	(x"93f20000", x"061e0000", x"44a0006c", x"65221800", x"07347453", x"36f6cc24", x"bb5dd99a", x"4484b662", x"be5d0000", x"ff4d0000", x"ed130057", x"67d02000", x"05dc6a7d", x"b16ebe19", x"15ae3bc7", x"34eab0f3"),
	(x"cbb10000", x"86600000", x"3c93006d", x"a3492000", x"e003288f", x"4f5bf3f9", x"172e27f5", x"7ec0cfd3", x"a3070000", x"d43f0000", x"a59e0057", x"c8b13800", x"201744b8", x"791701c9", x"940c3fee", x"2a9f8655"),
	(x"2b930000", x"394a0000", x"421d0072", x"b6ed0000", x"ad615743", x"8650d9c9", x"cdceb56b", x"51eac982", x"fca90000", x"e6110000", x"5ad9005c", x"99d70000", x"84523bca", x"487d50b0", x"cc07a3a3", x"80ae4e2a"),
	(x"73d00000", x"b9340000", x"3a2e0073", x"70863800", x"4a560b9f", x"fffde614", x"61bd4b04", x"6baeb033", x"e1f30000", x"cd630000", x"1254005c", x"36b61800", x"a199150f", x"8004ef60", x"4da5a78a", x"9edb788c"),
	(x"36c90000", x"12380000", x"0a900072", x"198c1800", x"88aa7986", x"4e296619", x"4c6cb142", x"4f9fff24", x"b9b00000", x"4d1d0000", x"6a67005d", x"f0dd2000", x"46ae49d3", x"f9a9d0bd", x"e1d659e5", x"a49f013d"),
	(x"6e8a0000", x"92460000", x"72a30073", x"dfe72000", x"6f9d255a", x"378459c4", x"e01f4f2d", x"75db8695", x"a4ea0000", x"666f0000", x"22ea005d", x"5fbc3800", x"63656716", x"31d06f6d", x"60745dcc", x"baea379b"),
	(x"0a1f0000", x"5bcb0000", x"8a1e0044", x"b3860000", x"01283651", x"a2673774", x"92728b63", x"f42251fd", x"d10a0000", x"eda30000", x"6b26006c", x"1e370000", x"fa943185", x"510c6bea", x"93a3bb17", x"6da573f8"),
	(x"525c0000", x"dbb50000", x"f22d0045", x"75ed3800", x"e61f6a8d", x"dbca08a9", x"3e01750c", x"ce66284c", x"cc500000", x"c6d10000", x"23ab006c", x"b1561800", x"df5f1f40", x"9975d43a", x"1201bf3e", x"73d0455e"),
	(x"17450000", x"70b90000", x"c2930044", x"1ce71800", x"24e31894", x"6a1e88a4", x"13d08f4a", x"ea57675b", x"94130000", x"46af0000", x"5b98006d", x"773d2000", x"3868439c", x"e0d8ebe7", x"be724151", x"49943cef"),
	(x"4f060000", x"f0c70000", x"baa00045", x"da8c2000", x"c3d44448", x"13b3b779", x"bfa37125", x"d0131eea", x"89490000", x"6ddd0000", x"1315006d", x"d85c3800", x"1da36d59", x"28a15437", x"3fd04578", x"57e10a49"),
	(x"af240000", x"4fed0000", x"c42e005a", x"cf280000", x"8eb63b84", x"dab89d49", x"6543e3bb", x"ff3918bb", x"d6e70000", x"5ff30000", x"ec520066", x"893a0000", x"b9e6122b", x"19cb054e", x"67dbd935", x"fdd0c236"),
	(x"f7670000", x"cf930000", x"bc1d005b", x"09433800", x"69816758", x"a315a294", x"c9301dd4", x"c57d610a", x"cbbd0000", x"74810000", x"a4df0066", x"265b1800", x"9c2d3cee", x"d1b2ba9e", x"e679dd1c", x"e3a5f490"),
	(x"b27e0000", x"649f0000", x"8ca3005a", x"60491800", x"ab7d1541", x"12c12299", x"e4e1e792", x"e14c2e1d", x"93fe0000", x"f4ff0000", x"dcec0067", x"e0302000", x"7b1a6032", x"a81f8543", x"4a0a2373", x"d9e18d21"),
	(x"ea3d0000", x"e4e10000", x"f490005b", x"a6222000", x"4c4a499d", x"6b6c1d44", x"489219fd", x"db0857ac", x"8ea40000", x"df8d0000", x"94610067", x"4f513800", x"5ed14ef7", x"60663a93", x"cba8275a", x"c794bb87"),
	(x"0df20000", x"e99b0000", x"0d6a004e", x"248b0000", x"425a15ff", x"eaa059d0", x"660ae941", x"6457e033", x"73dc0000", x"4bd50000", x"a2620078", x"f5940000", x"36781ffe", x"6114af73", x"90eab1ed", x"f6cb8b70"),
	(x"55b10000", x"69e50000", x"7559004f", x"e2e03800", x"a56d4923", x"930d660d", x"ca79172e", x"5e139982", x"6e860000", x"60a70000", x"eaef0078", x"5af51800", x"13b3313b", x"a96d10a3", x"1148b5c4", x"e8bebdd6"),
	(x"10a80000", x"c2e90000", x"45e7004e", x"8bea1800", x"67913b3a", x"22d9e600", x"e7a8ed68", x"7a22d695", x"36c50000", x"e0d90000", x"92dc0079", x"9c9e2000", x"f4846de7", x"d0c02f7e", x"bd3b4bab", x"d2fac467"),
	(x"48eb0000", x"42970000", x"3dd4004f", x"4d812000", x"80a667e6", x"5b74d9dd", x"4bdb1307", x"4066af24", x"2b9f0000", x"cbab0000", x"da510079", x"33ff3800", x"d14f4322", x"18b990ae", x"3c994f82", x"cc8ff2c1"),
	(x"a8c90000", x"fdbd0000", x"435a0050", x"58250000", x"cdc4182a", x"927ff3ed", x"913b8199", x"6f4ca975", x"74310000", x"f9850000", x"25160072", x"62990000", x"750a3c50", x"29d3c1d7", x"6492d3cf", x"66be3abe"),
	(x"f08a0000", x"7dc30000", x"3b690051", x"9e4e3800", x"2af344f6", x"ebd2cc30", x"3d487ff6", x"5508d0c4", x"696b0000", x"d2f70000", x"6d9b0072", x"cdf81800", x"50c11295", x"e1aa7e07", x"e530d7e6", x"78cb0c18"),
	(x"b5930000", x"d6cf0000", x"0bd70050", x"f7441800", x"e80f36ef", x"5a064c3d", x"109985b0", x"71399fd3", x"31280000", x"52890000", x"15a80073", x"0b932000", x"b7f64e49", x"980741da", x"49432989", x"428f75a9"),
	(x"edd00000", x"56b10000", x"73e40051", x"312f2000", x"0f386a33", x"23ab73e0", x"bcea7bdf", x"4b7de662", x"2c720000", x"79fb0000", x"5d250073", x"a4f23800", x"923d608c", x"507efe0a", x"c8e12da0", x"5cfa430f"),
	(x"82870000", x"445f0000", x"f5d1006a", x"48c80000", x"f07031cb", x"c3c9a613", x"3ae7fb0f", x"12322569", x"dac80000", x"36c00000", x"15ae0060", x"0bb10000", x"6b697976", x"248dd0a9", x"67c3ff89", x"b513679b"),
	(x"dac40000", x"c4210000", x"8de2006b", x"8ea33800", x"17476d17", x"ba6499ce", x"96940560", x"28765cd8", x"c7920000", x"1db20000", x"5d230060", x"a4d01800", x"4ea257b3", x"ecf46f79", x"e661fba0", x"ab66513d"),
	(x"9fdd0000", x"6f2d0000", x"bd5c006a", x"e7a91800", x"d5bb1f0e", x"0bb019c3", x"bb45ff26", x"0c4713cf", x"9fd10000", x"9dcc0000", x"25100061", x"62bb2000", x"a9950b6f", x"955950a4", x"4a1205cf", x"9122288c"),
	(x"c79e0000", x"ef530000", x"c56f006b", x"21c22000", x"328c43d2", x"721d261e", x"17360149", x"36036a7e", x"828b0000", x"b6be0000", x"6d9d0061", x"cdda3800", x"8c5e25aa", x"5d20ef74", x"cbb001e6", x"8f571e2a"),
	(x"27bc0000", x"50790000", x"bbe10074", x"34660000", x"7fee3c1e", x"bb160c2e", x"cdd693d7", x"19296c2f", x"dd250000", x"84900000", x"92da006a", x"9cbc0000", x"281b5ad8", x"6c4abe0d", x"93bb9dab", x"2566d655"),
	(x"7fff0000", x"d0070000", x"c3d20075", x"f20d3800", x"98d960c2", x"c2bb33f3", x"61a56db8", x"236d159e", x"c07f0000", x"afe20000", x"da57006a", x"33dd1800", x"0dd0741d", x"a43301dd", x"12199982", x"3b13e0f3"),
	(x"3ae60000", x"7b0b0000", x"f36c0074", x"9b071800", x"5a2512db", x"736fb3fe", x"4c7497fe", x"075c5a89", x"983c0000", x"2f9c0000", x"a264006b", x"f5b62000", x"eae728c1", x"dd9e3e00", x"be6a67ed", x"01579942"),
	(x"62a50000", x"fb750000", x"8b5f0075", x"5d6c2000", x"bd124e07", x"0ac28c23", x"e0076991", x"3d182338", x"85660000", x"04ee0000", x"eae9006b", x"5ad73800", x"cf2c0604", x"15e781d0", x"3fc863c4", x"1f22afe4"),
	(x"856a0000", x"f60f0000", x"72a50060", x"dfc50000", x"b3021265", x"8b0ec8b7", x"ce9f992d", x"824794a7", x"781e0000", x"90b60000", x"dcea0074", x"e0120000", x"a785570d", x"14951430", x"648af573", x"2e7d9f13"),
	(x"dd290000", x"76710000", x"0a960061", x"19ae3800", x"54354eb9", x"f2a3f76a", x"62ec6742", x"b803ed16", x"65440000", x"bbc40000", x"94670074", x"4f731800", x"824e79c8", x"dcecabe0", x"e528f15a", x"3008a9b5"),
	(x"98300000", x"dd7d0000", x"3a280060", x"70a41800", x"96c93ca0", x"43777767", x"4f3d9d04", x"9c32a201", x"3d070000", x"3bba0000", x"ec540075", x"89182000", x"65792514", x"a541943d", x"495b0f35", x"0a4cd004"),
	(x"c0730000", x"5d030000", x"421b0061", x"b6cf2000", x"71fe607c", x"3ada48ba", x"e34e636b", x"a676dbb0", x"205d0000", x"10c80000", x"a4d90075", x"26793800", x"40b20bd1", x"6d382bed", x"c8f90b1c", x"1439e6a2"),
	(x"20510000", x"e2290000", x"3c95007e", x"a36b0000", x"3c9c1fb0", x"f3d1628a", x"39aef1f5", x"895cdde1", x"7ff30000", x"22e60000", x"5b9e007e", x"771f0000", x"e4f774a3", x"5c527a94", x"90f29751", x"be082edd"),
	(x"78120000", x"62570000", x"44a6007f", x"65003800", x"dbab436c", x"8a7c5d57", x"95dd0f9a", x"b318a450", x"62a90000", x"09940000", x"1313007e", x"d87e1800", x"c13c5a66", x"942bc544", x"11509378", x"a07d187b"),
	(x"3d0b0000", x"c95b0000", x"7418007e", x"0c0a1800", x"19573175", x"3ba8dd5a", x"b80cf5dc", x"9729eb47", x"3aea0000", x"89ea0000", x"6b20007f", x"1e152000", x"260b06ba", x"ed86fa99", x"bd236d17", x"9a3961ca"),
	(x"65480000", x"49250000", x"0c2b007f", x"ca612000", x"fe606da9", x"4205e287", x"147f0bb3", x"ad6d92f6", x"27b00000", x"a2980000", x"23ad007f", x"b1743800", x"03c0287f", x"25ff4549", x"3c81693e", x"844c576c")
    ),(
	(x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000"),
	(x"e6280000", x"4c4b0000", x"a8550000", x"d3d002e0", x"d86130b8", x"98a7b0da", x"289506b4", x"d75a4897", x"f0c50000", x"59230000", x"45820000", x"e18d00c0", x"3b6d0631", x"c2ed5699", x"cbe0fe1c", x"56a7b19f"),
	(x"f0c50000", x"59230000", x"45820000", x"e18d00c0", x"3b6d0631", x"c2ed5699", x"cbe0fe1c", x"56a7b19f", x"16ed0000", x"15680000", x"edd70000", x"325d0220", x"e30c3689", x"5a4ae643", x"e375f8a8", x"81fdf908"),
	(x"16ed0000", x"15680000", x"edd70000", x"325d0220", x"e30c3689", x"5a4ae643", x"e375f8a8", x"81fdf908", x"e6280000", x"4c4b0000", x"a8550000", x"d3d002e0", x"d86130b8", x"98a7b0da", x"289506b4", x"d75a4897"),
	(x"b4310000", x"77330000", x"b15d0000", x"7fd004e0", x"78a26138", x"d116c35d", x"d256d489", x"4e6f74de", x"e3060000", x"bdc10000", x"87130000", x"bff20060", x"2eba0a1a", x"8db53751", x"73c5ab06", x"5bd61539"),
	(x"52190000", x"3b780000", x"19080000", x"ac000600", x"a0c35180", x"49b17387", x"fac3d23d", x"99353c49", x"13c30000", x"e4e20000", x"c2910000", x"5e7f00a0", x"15d70c2b", x"4f5861c8", x"b825551a", x"0d71a4a6"),
	(x"44f40000", x"2e100000", x"f4df0000", x"9e5d0420", x"43cf6709", x"13fb95c4", x"19b62a95", x"18c8c541", x"f5eb0000", x"a8a90000", x"6ac40000", x"8daf0240", x"cdb63c93", x"d7ffd112", x"90b053ae", x"da2bec31"),
	(x"a2dc0000", x"625b0000", x"5c8a0000", x"4d8d06c0", x"9bae57b1", x"8b5c251e", x"31232c21", x"cf928dd6", x"052e0000", x"f18a0000", x"2f460000", x"6c220280", x"f6db3aa2", x"1512878b", x"5b50adb2", x"8c8c5dae"),
	(x"e3060000", x"bdc10000", x"87130000", x"bff20060", x"2eba0a1a", x"8db53751", x"73c5ab06", x"5bd61539", x"57370000", x"caf20000", x"364e0000", x"c0220480", x"56186b22", x"5ca3f40c", x"a1937f8f", x"15b961e7"),
	(x"052e0000", x"f18a0000", x"2f460000", x"6c220280", x"f6db3aa2", x"1512878b", x"5b50adb2", x"8c8c5dae", x"a7f20000", x"93d10000", x"73cc0000", x"21af0440", x"6d756d13", x"9e4ea295", x"6a738193", x"431ed078"),
	(x"13c30000", x"e4e20000", x"c2910000", x"5e7f00a0", x"15d70c2b", x"4f5861c8", x"b825551a", x"0d71a4a6", x"41da0000", x"df9a0000", x"db990000", x"f27f06a0", x"b5145dab", x"06e9124f", x"42e68727", x"944498ef"),
	(x"f5eb0000", x"a8a90000", x"6ac40000", x"8daf0240", x"cdb63c93", x"d7ffd112", x"90b053ae", x"da2bec31", x"b11f0000", x"86b90000", x"9e1b0000", x"13f20660", x"8e795b9a", x"c40444d6", x"8906793b", x"c2e32970"),
	(x"57370000", x"caf20000", x"364e0000", x"c0220480", x"56186b22", x"5ca3f40c", x"a1937f8f", x"15b961e7", x"b4310000", x"77330000", x"b15d0000", x"7fd004e0", x"78a26138", x"d116c35d", x"d256d489", x"4e6f74de"),
	(x"b11f0000", x"86b90000", x"9e1b0000", x"13f20660", x"8e795b9a", x"c40444d6", x"8906793b", x"c2e32970", x"44f40000", x"2e100000", x"f4df0000", x"9e5d0420", x"43cf6709", x"13fb95c4", x"19b62a95", x"18c8c541"),
	(x"a7f20000", x"93d10000", x"73cc0000", x"21af0440", x"6d756d13", x"9e4ea295", x"6a738193", x"431ed078", x"a2dc0000", x"625b0000", x"5c8a0000", x"4d8d06c0", x"9bae57b1", x"8b5c251e", x"31232c21", x"cf928dd6"),
	(x"41da0000", x"df9a0000", x"db990000", x"f27f06a0", x"b5145dab", x"06e9124f", x"42e68727", x"944498ef", x"52190000", x"3b780000", x"19080000", x"ac000600", x"a0c35180", x"49b17387", x"fac3d23d", x"99353c49"),
	(x"02f20000", x"a2810000", x"873f0000", x"e36c7800", x"1e1d74ef", x"073d2bd6", x"c4c23237", x"7f32259e", x"badd0000", x"13ad0000", x"b7e70000", x"f7282800", x"df45144d", x"361ac33a", x"ea5a8d14", x"2a2c18f0"),
	(x"e4da0000", x"eeca0000", x"2f6a0000", x"30bc7ae0", x"c67c4457", x"9f9a9b0c", x"ec573483", x"a8686d09", x"4a180000", x"4a8e0000", x"f2650000", x"16a528c0", x"e428127c", x"f4f795a3", x"21ba7308", x"7c8ba96f"),
	(x"f2370000", x"fba20000", x"c2bd0000", x"02e178c0", x"257072de", x"c5d07d4f", x"0f22cc2b", x"29959401", x"ac300000", x"06c50000", x"5a300000", x"c5752a20", x"3c4922c4", x"6c502579", x"092f75bc", x"abd1e1f8"),
	(x"141f0000", x"b7e90000", x"6ae80000", x"d1317a20", x"fd114266", x"5d77cd95", x"27b7ca9f", x"fecfdc96", x"5cf50000", x"5fe60000", x"1fb20000", x"24f82ae0", x"072424f5", x"aebd73e0", x"c2cf8ba0", x"fd765067"),
	(x"b6c30000", x"d5b20000", x"36620000", x"9cbc7ce0", x"66bf15d7", x"d62be88b", x"1694e6be", x"315d5140", x"59db0000", x"ae6c0000", x"30f40000", x"48da2860", x"f1ff1e57", x"bbaff46b", x"999f2612", x"71fa0dc9"),
	(x"50eb0000", x"99f90000", x"9e370000", x"4f6c7e00", x"bede256f", x"4e8c5851", x"3e01e00a", x"e60719d7", x"a91e0000", x"f74f0000", x"75760000", x"a95728a0", x"ca921866", x"7942a2f2", x"527fd80e", x"275dbc56"),
	(x"46060000", x"8c910000", x"73e00000", x"7d317c20", x"5dd213e6", x"14c6be12", x"dd7418a2", x"67fae0df", x"4f360000", x"bb040000", x"dd230000", x"7a872a40", x"12f328de", x"e1e51228", x"7aeadeba", x"f007f4c1"),
	(x"a02e0000", x"c0da0000", x"dbb50000", x"aee17ec0", x"85b3235e", x"8c610ec8", x"f5e11e16", x"b0a0a848", x"bff30000", x"e2270000", x"98a10000", x"9b0a2a80", x"299e2eef", x"230844b1", x"b10a20a6", x"a6a0455e"),
	(x"e1f40000", x"1f400000", x"002c0000", x"5c9e7860", x"30a77ef5", x"8a881c87", x"b7079931", x"24e430a7", x"edea0000", x"d95f0000", x"81a90000", x"370a2c80", x"895d7f6f", x"6ab93736", x"4bc9f29b", x"3f957917"),
	(x"07dc0000", x"530b0000", x"a8790000", x"8f4e7a80", x"e8c64e4d", x"122fac5d", x"9f929f85", x"f3be7830", x"1d2f0000", x"807c0000", x"c42b0000", x"d6872c40", x"b230795e", x"a85461af", x"80290c87", x"6932c888"),
	(x"11310000", x"46630000", x"45ae0000", x"bd1378a0", x"0bca78c4", x"48654a1e", x"7ce7672d", x"72438138", x"fb070000", x"cc370000", x"6c7e0000", x"05572ea0", x"6a5149e6", x"30f3d175", x"a8bc0a33", x"be68801f"),
	(x"f7190000", x"0a280000", x"edfb0000", x"6ec37a40", x"d3ab487c", x"d0c2fac4", x"54726199", x"a519c9af", x"0bc20000", x"95140000", x"29fc0000", x"e4da2e60", x"513c4fd7", x"f21e87ec", x"635cf42f", x"e8cf3180"),
	(x"55c50000", x"68730000", x"b1710000", x"234e7c80", x"48051fcd", x"5b9edfda", x"65514db8", x"6a8b4479", x"0eec0000", x"649e0000", x"06ba0000", x"88f82ce0", x"a7e77575", x"e70c0067", x"380c599d", x"64436c2e"),
	(x"b3ed0000", x"24380000", x"19240000", x"f09e7e60", x"90642f75", x"c3396f00", x"4dc44b0c", x"bdd10cee", x"fe290000", x"3dbd0000", x"43380000", x"69752c20", x"9c8a7344", x"25e156fe", x"f3eca781", x"32e4ddb1"),
	(x"a5000000", x"31500000", x"f4f30000", x"c2c37c40", x"736819fc", x"99738943", x"aeb1b3a4", x"3c2cf5e6", x"18010000", x"71f60000", x"eb6d0000", x"baa52ec0", x"44eb43fc", x"bd46e624", x"db79a135", x"e5be9526"),
	(x"43280000", x"7d1b0000", x"5ca60000", x"11137ea0", x"ab092944", x"01d43999", x"8624b510", x"eb76bd71", x"e8c40000", x"28d50000", x"aeef0000", x"5b282e00", x"7f8645cd", x"7fabb0bd", x"10995f29", x"b31924b9"),
	(x"badd0000", x"13ad0000", x"b7e70000", x"f7282800", x"df45144d", x"361ac33a", x"ea5a8d14", x"2a2c18f0", x"b82f0000", x"b12c0000", x"30d80000", x"14445000", x"c15860a2", x"3127e8ec", x"2e98bf23", x"551e3d6e"),
	(x"5cf50000", x"5fe60000", x"1fb20000", x"24f82ae0", x"072424f5", x"aebd73e0", x"c2cf8ba0", x"fd765067", x"48ea0000", x"e80f0000", x"755a0000", x"f5c950c0", x"fa356693", x"f3cabe75", x"e578413f", x"03b98cf1"),
	(x"4a180000", x"4a8e0000", x"f2650000", x"16a528c0", x"e428127c", x"f4f795a3", x"21ba7308", x"7c8ba96f", x"aec20000", x"a4440000", x"dd0f0000", x"26195220", x"2254562b", x"6b6d0eaf", x"cded478b", x"d4e3c466"),
	(x"ac300000", x"06c50000", x"5a300000", x"c5752a20", x"3c4922c4", x"6c502579", x"092f75bc", x"abd1e1f8", x"5e070000", x"fd670000", x"988d0000", x"c79452e0", x"1939501a", x"a9805836", x"060db997", x"824475f9"),
	(x"0eec0000", x"649e0000", x"06ba0000", x"88f82ce0", x"a7e77575", x"e70c0067", x"380c599d", x"64436c2e", x"5b290000", x"0ced0000", x"b7cb0000", x"abb65060", x"efe26ab8", x"bc92dfbd", x"5d5d1425", x"0ec82857"),
	(x"e8c40000", x"28d50000", x"aeef0000", x"5b282e00", x"7f8645cd", x"7fabb0bd", x"10995f29", x"b31924b9", x"abec0000", x"55ce0000", x"f2490000", x"4a3b50a0", x"d48f6c89", x"7e7f8924", x"96bdea39", x"586f99c8"),
	(x"fe290000", x"3dbd0000", x"43380000", x"69752c20", x"9c8a7344", x"25e156fe", x"f3eca781", x"32e4ddb1", x"4dc40000", x"19850000", x"5a1c0000", x"99eb5240", x"0cee5c31", x"e6d839fe", x"be28ec8d", x"8f35d15f"),
	(x"18010000", x"71f60000", x"eb6d0000", x"baa52ec0", x"44eb43fc", x"bd46e624", x"db79a135", x"e5be9526", x"bd010000", x"40a60000", x"1f9e0000", x"78665280", x"37835a00", x"24356f67", x"75c81291", x"d99260c0"),
	(x"59db0000", x"ae6c0000", x"30f40000", x"48da2860", x"f1ff1e57", x"bbaff46b", x"999f2612", x"71fa0dc9", x"ef180000", x"7bde0000", x"06960000", x"d4665480", x"97400b80", x"6d841ce0", x"8f0bc0ac", x"40a75c89"),
	(x"bff30000", x"e2270000", x"98a10000", x"9b0a2a80", x"299e2eef", x"230844b1", x"b10a20a6", x"a6a0455e", x"1fdd0000", x"22fd0000", x"43140000", x"35eb5440", x"ac2d0db1", x"af694a79", x"44eb3eb0", x"1600ed16"),
	(x"a91e0000", x"f74f0000", x"75760000", x"a95728a0", x"ca921866", x"7942a2f2", x"527fd80e", x"275dbc56", x"f9f50000", x"6eb60000", x"eb410000", x"e63b56a0", x"744c3d09", x"37cefaa3", x"6c7e3804", x"c15aa581"),
	(x"4f360000", x"bb040000", x"dd230000", x"7a872a40", x"12f328de", x"e1e51228", x"7aeadeba", x"f007f4c1", x"09300000", x"37950000", x"aec30000", x"07b65660", x"4f213b38", x"f523ac3a", x"a79ec618", x"97fd141e"),
	(x"edea0000", x"d95f0000", x"81a90000", x"370a2c80", x"895d7f6f", x"6ab93736", x"4bc9f29b", x"3f957917", x"0c1e0000", x"c61f0000", x"81850000", x"6b9454e0", x"b9fa019a", x"e0312bb1", x"fcce6baa", x"1b7149b0"),
	(x"0bc20000", x"95140000", x"29fc0000", x"e4da2e60", x"513c4fd7", x"f21e87ec", x"635cf42f", x"e8cf3180", x"fcdb0000", x"9f3c0000", x"c4070000", x"8a195420", x"829707ab", x"22dc7d28", x"372e95b6", x"4dd6f82f"),
	(x"1d2f0000", x"807c0000", x"c42b0000", x"d6872c40", x"b230795e", x"a85461af", x"80290c87", x"6932c888", x"1af30000", x"d3770000", x"6c520000", x"59c956c0", x"5af63713", x"ba7bcdf2", x"1fbb9302", x"9a8cb0b8"),
	(x"fb070000", x"cc370000", x"6c7e0000", x"05572ea0", x"6a5149e6", x"30f3d175", x"a8bc0a33", x"be68801f", x"ea360000", x"8a540000", x"29d00000", x"b8445600", x"619b3122", x"78969b6b", x"d45b6d1e", x"cc2b0127"),
	(x"b82f0000", x"b12c0000", x"30d80000", x"14445000", x"c15860a2", x"3127e8ec", x"2e98bf23", x"551e3d6e", x"02f20000", x"a2810000", x"873f0000", x"e36c7800", x"1e1d74ef", x"073d2bd6", x"c4c23237", x"7f32259e"),
	(x"5e070000", x"fd670000", x"988d0000", x"c79452e0", x"1939501a", x"a9805836", x"060db997", x"824475f9", x"f2370000", x"fba20000", x"c2bd0000", x"02e178c0", x"257072de", x"c5d07d4f", x"0f22cc2b", x"29959401"),
	(x"48ea0000", x"e80f0000", x"755a0000", x"f5c950c0", x"fa356693", x"f3cabe75", x"e578413f", x"03b98cf1", x"141f0000", x"b7e90000", x"6ae80000", x"d1317a20", x"fd114266", x"5d77cd95", x"27b7ca9f", x"fecfdc96"),
	(x"aec20000", x"a4440000", x"dd0f0000", x"26195220", x"2254562b", x"6b6d0eaf", x"cded478b", x"d4e3c466", x"e4da0000", x"eeca0000", x"2f6a0000", x"30bc7ae0", x"c67c4457", x"9f9a9b0c", x"ec573483", x"a8686d09"),
	(x"0c1e0000", x"c61f0000", x"81850000", x"6b9454e0", x"b9fa019a", x"e0312bb1", x"fcce6baa", x"1b7149b0", x"e1f40000", x"1f400000", x"002c0000", x"5c9e7860", x"30a77ef5", x"8a881c87", x"b7079931", x"24e430a7"),
	(x"ea360000", x"8a540000", x"29d00000", x"b8445600", x"619b3122", x"78969b6b", x"d45b6d1e", x"cc2b0127", x"11310000", x"46630000", x"45ae0000", x"bd1378a0", x"0bca78c4", x"48654a1e", x"7ce7672d", x"72438138"),
	(x"fcdb0000", x"9f3c0000", x"c4070000", x"8a195420", x"829707ab", x"22dc7d28", x"372e95b6", x"4dd6f82f", x"f7190000", x"0a280000", x"edfb0000", x"6ec37a40", x"d3ab487c", x"d0c2fac4", x"54726199", x"a519c9af"),
	(x"1af30000", x"d3770000", x"6c520000", x"59c956c0", x"5af63713", x"ba7bcdf2", x"1fbb9302", x"9a8cb0b8", x"07dc0000", x"530b0000", x"a8790000", x"8f4e7a80", x"e8c64e4d", x"122fac5d", x"9f929f85", x"f3be7830"),
	(x"5b290000", x"0ced0000", x"b7cb0000", x"abb65060", x"efe26ab8", x"bc92dfbd", x"5d5d1425", x"0ec82857", x"55c50000", x"68730000", x"b1710000", x"234e7c80", x"48051fcd", x"5b9edfda", x"65514db8", x"6a8b4479"),
	(x"bd010000", x"40a60000", x"1f9e0000", x"78665280", x"37835a00", x"24356f67", x"75c81291", x"d99260c0", x"a5000000", x"31500000", x"f4f30000", x"c2c37c40", x"736819fc", x"99738943", x"aeb1b3a4", x"3c2cf5e6"),
	(x"abec0000", x"55ce0000", x"f2490000", x"4a3b50a0", x"d48f6c89", x"7e7f8924", x"96bdea39", x"586f99c8", x"43280000", x"7d1b0000", x"5ca60000", x"11137ea0", x"ab092944", x"01d43999", x"8624b510", x"eb76bd71"),
	(x"4dc40000", x"19850000", x"5a1c0000", x"99eb5240", x"0cee5c31", x"e6d839fe", x"be28ec8d", x"8f35d15f", x"b3ed0000", x"24380000", x"19240000", x"f09e7e60", x"90642f75", x"c3396f00", x"4dc44b0c", x"bdd10cee"),
	(x"ef180000", x"7bde0000", x"06960000", x"d4665480", x"97400b80", x"6d841ce0", x"8f0bc0ac", x"40a75c89", x"b6c30000", x"d5b20000", x"36620000", x"9cbc7ce0", x"66bf15d7", x"d62be88b", x"1694e6be", x"315d5140"),
	(x"09300000", x"37950000", x"aec30000", x"07b65660", x"4f213b38", x"f523ac3a", x"a79ec618", x"97fd141e", x"46060000", x"8c910000", x"73e00000", x"7d317c20", x"5dd213e6", x"14c6be12", x"dd7418a2", x"67fae0df"),
	(x"1fdd0000", x"22fd0000", x"43140000", x"35eb5440", x"ac2d0db1", x"af694a79", x"44eb3eb0", x"1600ed16", x"a02e0000", x"c0da0000", x"dbb50000", x"aee17ec0", x"85b3235e", x"8c610ec8", x"f5e11e16", x"b0a0a848"),
	(x"f9f50000", x"6eb60000", x"eb410000", x"e63b56a0", x"744c3d09", x"37cefaa3", x"6c7e3804", x"c15aa581", x"50eb0000", x"99f90000", x"9e370000", x"4f6c7e00", x"bede256f", x"4e8c5851", x"3e01e00a", x"e60719d7"),
	(x"1e6c0000", x"c4420000", x"8a2e0000", x"bcb6b800", x"2c4413b6", x"8bfdd3da", x"6a0c1bc8", x"b99dc2eb", x"92560000", x"1eda0000", x"ea510000", x"e8b13000", x"a93556a5", x"ebfb6199", x"b15c2254", x"33c5244f"),
	(x"f8440000", x"88090000", x"227b0000", x"6f66bae0", x"f425230e", x"135a6300", x"42991d7c", x"6ec78a7c", x"62930000", x"47f90000", x"afd30000", x"093c30c0", x"92585094", x"29163700", x"7abcdc48", x"656295d0"),
	(x"eea90000", x"9d610000", x"cfac0000", x"5d3bb8c0", x"17291587", x"49108543", x"a1ece5d4", x"ef3a7374", x"84bb0000", x"0bb20000", x"07860000", x"daec3220", x"4a39602c", x"b1b187da", x"5229dafc", x"b238dd47"),
	(x"08810000", x"d12a0000", x"67f90000", x"8eebba20", x"cf48253f", x"d1b73599", x"8979e360", x"38603be3", x"747e0000", x"52910000", x"42040000", x"3b6132e0", x"7154661d", x"735cd143", x"99c924e0", x"e49f6cd8"),
	(x"aa5d0000", x"b3710000", x"3b730000", x"c366bce0", x"54e6728e", x"5aeb1087", x"b85acf41", x"f7f2b635", x"71500000", x"a31b0000", x"6d420000", x"57433060", x"878f5cbf", x"664e56c8", x"c2998952", x"68133176"),
	(x"4c750000", x"ff3a0000", x"93260000", x"10b6be00", x"8c874236", x"c24ca05d", x"90cfc9f5", x"20a8fea2", x"81950000", x"fa380000", x"28c00000", x"b6ce30a0", x"bce25a8e", x"a4a30051", x"0979774e", x"3eb480e9"),
	(x"5a980000", x"ea520000", x"7ef10000", x"22ebbc20", x"6f8b74bf", x"9806461e", x"73ba315d", x"a15507aa", x"67bd0000", x"b6730000", x"80950000", x"651e3240", x"64836a36", x"3c04b08b", x"21ec71fa", x"e9eec87e"),
	(x"bcb00000", x"a6190000", x"d6a40000", x"f13bbec0", x"b7ea4407", x"00a1f6c4", x"5b2f37e9", x"760f4f3d", x"97780000", x"ef500000", x"c5170000", x"84933280", x"5fee6c07", x"fee9e612", x"ea0c8fe6", x"bf4979e1"),
	(x"fd6a0000", x"79830000", x"0d3d0000", x"0344b860", x"02fe19ac", x"0648e48b", x"19c9b0ce", x"e24bd7d2", x"c5610000", x"d4280000", x"dc1f0000", x"28933480", x"ff2d3d87", x"b7589595", x"10cf5ddb", x"267c45a8"),
	(x"1b420000", x"35c80000", x"a5680000", x"d094ba80", x"da9f2914", x"9eef5451", x"315cb67a", x"35119f45", x"35a40000", x"8d0b0000", x"999d0000", x"c91e3440", x"c4403bb6", x"75b5c30c", x"db2fa3c7", x"70dbf437"),
	(x"0daf0000", x"20a00000", x"48bf0000", x"e2c9b8a0", x"39931f9d", x"c4a5b212", x"d2294ed2", x"b4ec664d", x"d38c0000", x"c1400000", x"31c80000", x"1ace36a0", x"1c210b0e", x"ed1273d6", x"f3baa573", x"a781bca0"),
	(x"eb870000", x"6ceb0000", x"e0ea0000", x"3119ba40", x"e1f22f25", x"5c0202c8", x"fabc4866", x"63b62eda", x"23490000", x"98630000", x"744a0000", x"fb433660", x"274c0d3f", x"2fff254f", x"385a5b6f", x"f1260d3f"),
	(x"495b0000", x"0eb00000", x"bc600000", x"7c94bc80", x"7a5c7894", x"d75e27d6", x"cb9f6447", x"ac24a30c", x"26670000", x"69e90000", x"5b0c0000", x"976134e0", x"d197379d", x"3aeda2c4", x"630af6dd", x"7daa5091"),
	(x"af730000", x"42fb0000", x"14350000", x"af44be60", x"a23d482c", x"4ff9970c", x"e30a62f3", x"7b7eeb9b", x"d6a20000", x"30ca0000", x"1e8e0000", x"76ec3420", x"eafa31ac", x"f800f45d", x"a8ea08c1", x"2b0de10e"),
	(x"b99e0000", x"57930000", x"f9e20000", x"9d19bc40", x"41317ea5", x"15b3714f", x"007f9a5b", x"fa831293", x"308a0000", x"7c810000", x"b6db0000", x"a53c36c0", x"329b0114", x"60a74487", x"807f0e75", x"fc57a999"),
	(x"5fb60000", x"1bd80000", x"51b70000", x"4ec9bea0", x"99504e1d", x"8d14c195", x"28ea9cef", x"2dd95a04", x"c04f0000", x"25a20000", x"f3590000", x"44b13600", x"09f60725", x"a24a121e", x"4b9ff069", x"aaf01806"),
	(x"1c9e0000", x"66c30000", x"0d110000", x"5fdac000", x"32596759", x"8cc0f80c", x"aece29ff", x"c6afe775", x"288b0000", x"0d770000", x"5db60000", x"1f991800", x"767042e8", x"dde1a2a3", x"5b06af40", x"19e93cbf"),
	(x"fab60000", x"2a880000", x"a5440000", x"8c0ac2e0", x"ea3857e1", x"146748d6", x"865b2f4b", x"11f5afe2", x"d84e0000", x"54540000", x"18340000", x"fe1418c0", x"4d1d44d9", x"1f0cf43a", x"90e6515c", x"4f4e8d20"),
	(x"ec5b0000", x"3fe00000", x"48930000", x"be57c0c0", x"09346168", x"4e2dae95", x"652ed7e3", x"900856ea", x"3e660000", x"181f0000", x"b0610000", x"2dc41a20", x"957c7461", x"87ab44e0", x"b87357e8", x"9814c5b7"),
	(x"0a730000", x"73ab0000", x"e0c60000", x"6d87c220", x"d15551d0", x"d68a1e4f", x"4dbbd157", x"47521e7d", x"cea30000", x"413c0000", x"f5e30000", x"cc491ae0", x"ae117250", x"45461279", x"7393a9f4", x"ceb37428"),
	(x"a8af0000", x"11f00000", x"bc4c0000", x"200ac4e0", x"4afb0661", x"5dd63b51", x"7c98fd76", x"88c093ab", x"cb8d0000", x"b0b60000", x"daa50000", x"a06b1860", x"58ca48f2", x"505495f2", x"28c30446", x"423f2986"),
	(x"4e870000", x"5dbb0000", x"14190000", x"f3dac600", x"929a36d9", x"c5718b8b", x"540dfbc2", x"5f9adb3c", x"3b480000", x"e9950000", x"9f270000", x"41e618a0", x"63a74ec3", x"92b9c36b", x"e323fa5a", x"14989819"),
	(x"586a0000", x"48d30000", x"f9ce0000", x"c187c420", x"71960050", x"9f3b6dc8", x"b778036a", x"de672234", x"dd600000", x"a5de0000", x"37720000", x"92361a40", x"bbc67e7b", x"0a1e73b1", x"cbb6fcee", x"c3c2d08e"),
	(x"be420000", x"04980000", x"519b0000", x"1257c6c0", x"a9f730e8", x"079cdd12", x"9fed05de", x"093d6aa3", x"2da50000", x"fcfd0000", x"72f00000", x"73bb1a80", x"80ab784a", x"c8f32528", x"005602f2", x"95656111"),
	(x"ff980000", x"db020000", x"8a020000", x"e028c060", x"1ce36d43", x"0175cf5d", x"dd0b82f9", x"9d79f24c", x"7fbc0000", x"c7850000", x"6bf80000", x"dfbb1c80", x"206829ca", x"814256af", x"fa95d0cf", x"0c505d58"),
	(x"19b00000", x"97490000", x"22570000", x"33f8c280", x"c4825dfb", x"99d27f87", x"f59e844d", x"4a23badb", x"8f790000", x"9ea60000", x"2e7a0000", x"3e361c40", x"1b052ffb", x"43af0036", x"31752ed3", x"5af7ecc7"),
	(x"0f5d0000", x"82210000", x"cf800000", x"01a5c0a0", x"278e6b72", x"c39899c4", x"16eb7ce5", x"cbde43d3", x"69510000", x"d2ed0000", x"862f0000", x"ede61ea0", x"c3641f43", x"db08b0ec", x"19e02867", x"8dada450"),
	(x"e9750000", x"ce6a0000", x"67d50000", x"d275c240", x"ffef5bca", x"5b3f291e", x"3e7e7a51", x"1c840b44", x"99940000", x"8bce0000", x"c3ad0000", x"0c6b1e60", x"f8091972", x"19e5e675", x"d200d67b", x"db0a15cf"),
	(x"4ba90000", x"ac310000", x"3b5f0000", x"9ff8c480", x"64410c7b", x"d0630c00", x"0f5d5670", x"d3168692", x"9cba0000", x"7a440000", x"eceb0000", x"60491ce0", x"0ed223d0", x"0cf761fe", x"89507bc9", x"57864861"),
	(x"ad810000", x"e07a0000", x"930a0000", x"4c28c660", x"bc203cc3", x"48c4bcda", x"27c850c4", x"044cce05", x"6c7f0000", x"23670000", x"a9690000", x"81c41c20", x"35bf25e1", x"ce1a3767", x"42b085d5", x"0121f9fe"),
	(x"bb6c0000", x"f5120000", x"7edd0000", x"7e75c440", x"5f2c0a4a", x"128e5a99", x"c4bda86c", x"85b1370d", x"8a570000", x"6f2c0000", x"013c0000", x"52141ec0", x"edde1559", x"56bd87bd", x"6a258361", x"d67bb169"),
	(x"5d440000", x"b9590000", x"d6880000", x"ada5c6a0", x"874d3af2", x"8a29ea43", x"ec28aed8", x"52eb7f9a", x"7a920000", x"360f0000", x"44be0000", x"b3991e00", x"d6b31368", x"9450d124", x"a1c57d7d", x"80dc00f6"),
	(x"a4b10000", x"d7ef0000", x"3dc90000", x"4b9e9000", x"f30107fb", x"bde710e0", x"805696dc", x"93b1da1b", x"2a790000", x"aff60000", x"da890000", x"fcf56000", x"686d3607", x"dadc8975", x"9fc49d77", x"66db1921"),
	(x"42990000", x"9ba40000", x"959c0000", x"984e92e0", x"2b603743", x"2540a03a", x"a8c39068", x"44eb928c", x"dabc0000", x"f6d50000", x"9f0b0000", x"1d7860c0", x"53003036", x"1831dfec", x"5424636b", x"307ca8be"),
	(x"54740000", x"8ecc0000", x"784b0000", x"aa1390c0", x"c86c01ca", x"7f0a4679", x"4bb668c0", x"c5166b84", x"3c940000", x"ba9e0000", x"375e0000", x"cea86220", x"8b61008e", x"80966f36", x"7cb165df", x"e726e029"),
	(x"b25c0000", x"c2870000", x"d01e0000", x"79c39220", x"100d3172", x"e7adf6a3", x"63236e74", x"124c2313", x"cc510000", x"e3bd0000", x"72dc0000", x"2f2562e0", x"b00c06bf", x"427b39af", x"b7519bc3", x"b18151b6"),
	(x"10800000", x"a0dc0000", x"8c940000", x"344e94e0", x"8ba366c3", x"6cf1d3bd", x"52004255", x"dddeaec5", x"c97f0000", x"12370000", x"5d9a0000", x"43076060", x"46d73c1d", x"5769be24", x"ec013671", x"3d0d0c18"),
	(x"f6a80000", x"ec970000", x"24c10000", x"e79e9600", x"53c2567b", x"f4566367", x"7a9544e1", x"0a84e652", x"39ba0000", x"4b140000", x"18180000", x"a28a60a0", x"7dba3a2c", x"9584e8bd", x"27e1c86d", x"6baabd87"),
	(x"e0450000", x"f9ff0000", x"c9160000", x"d5c39420", x"b0ce60f2", x"ae1c8524", x"99e0bc49", x"8b791f5a", x"df920000", x"075f0000", x"b04d0000", x"715a6240", x"a5db0a94", x"0d235867", x"0f74ced9", x"bcf0f510"),
	(x"066d0000", x"b5b40000", x"61430000", x"061396c0", x"68af504a", x"36bb35fe", x"b175bafd", x"5c2357cd", x"2f570000", x"5e7c0000", x"f5cf0000", x"90d76280", x"9eb60ca5", x"cfce0efe", x"c49430c5", x"ea57448f"),
	(x"47b70000", x"6a2e0000", x"bada0000", x"f46c9060", x"ddbb0de1", x"305227b1", x"f3933dda", x"c867cf22", x"7d4e0000", x"65040000", x"ecc70000", x"3cd76480", x"3e755d25", x"867f7d79", x"3e57e2f8", x"736278c6"),
	(x"a19f0000", x"26650000", x"128f0000", x"27bc9280", x"05da3d59", x"a8f5976b", x"db063b6e", x"1f3d87b5", x"8d8b0000", x"3c270000", x"a9450000", x"dd5a6440", x"05185b14", x"44922be0", x"f5b71ce4", x"25c5c959"),
	(x"b7720000", x"330d0000", x"ff580000", x"15e190a0", x"e6d60bd0", x"f2bf7128", x"3873c3c6", x"9ec07ebd", x"6ba30000", x"706c0000", x"01100000", x"0e8a66a0", x"dd796bac", x"dc359b3a", x"dd221a50", x"f29f81ce"),
	(x"515a0000", x"7f460000", x"570d0000", x"c6319240", x"3eb73b68", x"6a18c1f2", x"10e6c572", x"499a362a", x"9b660000", x"294f0000", x"44920000", x"ef076660", x"e6146d9d", x"1ed8cda3", x"16c2e44c", x"a4383051"),
	(x"f3860000", x"1d1d0000", x"0b870000", x"8bbc9480", x"a5196cd9", x"e144e4ec", x"21c5e953", x"8608bbfc", x"9e480000", x"d8c50000", x"6bd40000", x"832564e0", x"10cf573f", x"0bca4a28", x"4d9249fe", x"28b46dff"),
	(x"15ae0000", x"51560000", x"a3d20000", x"586c9660", x"7d785c61", x"79e35436", x"0950efe7", x"5152f36b", x"6e8d0000", x"81e60000", x"2e560000", x"62a86420", x"2ba2510e", x"c9271cb1", x"8672b7e2", x"7e13dc60"),
	(x"03430000", x"443e0000", x"4e050000", x"6a319440", x"9e746ae8", x"23a9b275", x"ea25174f", x"d0af0a63", x"88a50000", x"cdad0000", x"86030000", x"b17866c0", x"f3c361b6", x"5180ac6b", x"aee7b156", x"a94994f7"),
	(x"e56b0000", x"08750000", x"e6500000", x"b9e196a0", x"46155a50", x"bb0e02af", x"c2b011fb", x"07f542f4", x"78600000", x"948e0000", x"c3810000", x"50f56600", x"c8ae6787", x"936dfaf2", x"65074f4a", x"ffee2568"),
	(x"a6430000", x"756e0000", x"baf60000", x"a8f2e800", x"ed1c7314", x"bada3b36", x"4494a4eb", x"ec83ff85", x"90a40000", x"bc5b0000", x"6d6e0000", x"0bdd4800", x"b728224a", x"ecc64a4f", x"759e1063", x"4cf701d1"),
	(x"406b0000", x"39250000", x"12a30000", x"7b22eae0", x"357d43ac", x"227d8bec", x"6c01a25f", x"3bd9b712", x"60610000", x"e5780000", x"28ec0000", x"ea5048c0", x"8c45247b", x"2e2b1cd6", x"be7eee7f", x"1a50b04e"),
	(x"56860000", x"2c4d0000", x"ff740000", x"497fe8c0", x"d6717525", x"78376daf", x"8f745af7", x"ba244e1a", x"86490000", x"a9330000", x"80b90000", x"39804a20", x"542414c3", x"b68cac0c", x"96ebe8cb", x"cd0af8d9"),
	(x"b0ae0000", x"60060000", x"57210000", x"9aafea20", x"0e10459d", x"e090dd75", x"a7e15c43", x"6d7e068d", x"768c0000", x"f0100000", x"c53b0000", x"d80d4ae0", x"6f4912f2", x"7461fa95", x"5d0b16d7", x"9bad4946"),
	(x"12720000", x"025d0000", x"0bab0000", x"d722ece0", x"95be122c", x"6bccf86b", x"96c27062", x"a2ec8b5b", x"73a20000", x"019a0000", x"ea7d0000", x"b42f4860", x"99922850", x"61737d1e", x"065bbb65", x"172114e8"),
	(x"f45a0000", x"4e160000", x"a3fe0000", x"04f2ee00", x"4ddf2294", x"f36b48b1", x"be5776d6", x"75b6c3cc", x"83670000", x"58b90000", x"afff0000", x"55a248a0", x"a2ff2e61", x"a39e2b87", x"cdbb4579", x"4186a577"),
	(x"e2b70000", x"5b7e0000", x"4e290000", x"36afec20", x"aed3141d", x"a921aef2", x"5d228e7e", x"f44b3ac4", x"654f0000", x"14f20000", x"07aa0000", x"86724a40", x"7a9e1ed9", x"3b399b5d", x"e52e43cd", x"96dcede0"),
	(x"049f0000", x"17350000", x"e67c0000", x"e57feec0", x"76b224a5", x"31861e28", x"75b788ca", x"23117253", x"958a0000", x"4dd10000", x"42280000", x"67ff4a80", x"41f318e8", x"f9d4cdc4", x"2ecebdd1", x"c07b5c7f"),
	(x"45450000", x"c8af0000", x"3de50000", x"1700e860", x"c3a6790e", x"376f0c67", x"37510fed", x"b755eabc", x"c7930000", x"76a90000", x"5b200000", x"cbff4c80", x"e1304968", x"b065be43", x"d40d6fec", x"594e6036"),
	(x"a36d0000", x"84e40000", x"95b00000", x"c4d0ea80", x"1bc749b6", x"afc8bcbd", x"1fc40959", x"600fa22b", x"37560000", x"2f8a0000", x"1ea20000", x"2a724c40", x"da5d4f59", x"7288e8da", x"1fed91f0", x"0fe9d1a9"),
	(x"b5800000", x"918c0000", x"78670000", x"f68de8a0", x"f8cb7f3f", x"f5825afe", x"fcb1f1f1", x"e1f25b23", x"d17e0000", x"63c10000", x"b6f70000", x"f9a24ea0", x"023c7fe1", x"ea2f5800", x"37789744", x"d8b3993e"),
	(x"53a80000", x"ddc70000", x"d0320000", x"255dea40", x"20aa4f87", x"6d25ea24", x"d424f745", x"36a813b4", x"21bb0000", x"3ae20000", x"f3750000", x"182f4e60", x"395179d0", x"28c20e99", x"fc986958", x"8e1428a1"),
	(x"f1740000", x"bf9c0000", x"8cb80000", x"68d0ec80", x"bb041836", x"e679cf3a", x"e507db64", x"f93a9e62", x"24950000", x"cb680000", x"dc330000", x"740d4ce0", x"cf8a4372", x"3dd08912", x"a7c8c4ea", x"0298750f"),
	(x"175c0000", x"f3d70000", x"24ed0000", x"bb00ee60", x"6365288e", x"7ede7fe0", x"cd92ddd0", x"2e60d6f5", x"d4500000", x"924b0000", x"99b10000", x"95804c20", x"f4e74543", x"ff3ddf8b", x"6c283af6", x"543fc490"),
	(x"01b10000", x"e6bf0000", x"c93a0000", x"895dec40", x"80691e07", x"249499a3", x"2ee72578", x"af9d2ffd", x"32780000", x"de000000", x"31e40000", x"46504ec0", x"2c8675fb", x"679a6f51", x"44bd3c42", x"83658c07"),
	(x"e7990000", x"aaf40000", x"616f0000", x"5a8deea0", x"58082ebf", x"bc332979", x"067223cc", x"78c7676a", x"c2bd0000", x"87230000", x"74660000", x"a7dd4e00", x"17eb73ca", x"a57739c8", x"8f5dc25e", x"d5c23d98"),
	(x"92560000", x"1eda0000", x"ea510000", x"e8b13000", x"a93556a5", x"ebfb6199", x"b15c2254", x"33c5244f", x"8c3a0000", x"da980000", x"607f0000", x"54078800", x"85714513", x"6006b243", x"db50399c", x"8a58e6a4"),
	(x"747e0000", x"52910000", x"42040000", x"3b6132e0", x"7154661d", x"735cd143", x"99c924e0", x"e49f6cd8", x"7cff0000", x"83bb0000", x"25fd0000", x"b58a88c0", x"be1c4322", x"a2ebe4da", x"10b0c780", x"dcff573b"),
	(x"62930000", x"47f90000", x"afd30000", x"093c30c0", x"92585094", x"29163700", x"7abcdc48", x"656295d0", x"9ad70000", x"cff00000", x"8da80000", x"665a8a20", x"667d739a", x"3a4c5400", x"3825c134", x"0ba51fac"),
	(x"84bb0000", x"0bb20000", x"07860000", x"daec3220", x"4a39602c", x"b1b187da", x"5229dafc", x"b238dd47", x"6a120000", x"96d30000", x"c82a0000", x"87d78ae0", x"5d1075ab", x"f8a10299", x"f3c53f28", x"5d02ae33"),
	(x"26670000", x"69e90000", x"5b0c0000", x"976134e0", x"d197379d", x"3aeda2c4", x"630af6dd", x"7daa5091", x"6f3c0000", x"67590000", x"e76c0000", x"ebf58860", x"abcb4f09", x"edb38512", x"a895929a", x"d18ef39d"),
	(x"c04f0000", x"25a20000", x"f3590000", x"44b13600", x"09f60725", x"a24a121e", x"4b9ff069", x"aaf01806", x"9ff90000", x"3e7a0000", x"a2ee0000", x"0a7888a0", x"90a64938", x"2f5ed38b", x"63756c86", x"87294202"),
	(x"d6a20000", x"30ca0000", x"1e8e0000", x"76ec3420", x"eafa31ac", x"f800f45d", x"a8ea08c1", x"2b0de10e", x"79d10000", x"72310000", x"0abb0000", x"d9a88a40", x"48c77980", x"b7f96351", x"4be06a32", x"50730a95"),
	(x"308a0000", x"7c810000", x"b6db0000", x"a53c36c0", x"329b0114", x"60a74487", x"807f0e75", x"fc57a999", x"89140000", x"2b120000", x"4f390000", x"38258a80", x"73aa7fb1", x"751435c8", x"8000942e", x"06d4bb0a"),
	(x"71500000", x"a31b0000", x"6d420000", x"57433060", x"878f5cbf", x"664e56c8", x"c2998952", x"68133176", x"db0d0000", x"106a0000", x"56310000", x"94258c80", x"d3692e31", x"3ca5464f", x"7ac34613", x"9fe18743"),
	(x"97780000", x"ef500000", x"c5170000", x"84933280", x"5fee6c07", x"fee9e612", x"ea0c8fe6", x"bf4979e1", x"2bc80000", x"49490000", x"13b30000", x"75a88c40", x"e8042800", x"fe4810d6", x"b123b80f", x"c94636dc"),
	(x"81950000", x"fa380000", x"28c00000", x"b6ce30a0", x"bce25a8e", x"a4a30051", x"0979774e", x"3eb480e9", x"cde00000", x"05020000", x"bbe60000", x"a6788ea0", x"306518b8", x"66efa00c", x"99b6bebb", x"1e1c7e4b"),
	(x"67bd0000", x"b6730000", x"80950000", x"651e3240", x"64836a36", x"3c04b08b", x"21ec71fa", x"e9eec87e", x"3d250000", x"5c210000", x"fe640000", x"47f58e60", x"0b081e89", x"a402f695", x"525640a7", x"48bbcfd4"),
	(x"c5610000", x"d4280000", x"dc1f0000", x"28933480", x"ff2d3d87", x"b7589595", x"10cf5ddb", x"267c45a8", x"380b0000", x"adab0000", x"d1220000", x"2bd78ce0", x"fdd3242b", x"b110711e", x"0906ed15", x"c437927a"),
	(x"23490000", x"98630000", x"744a0000", x"fb433660", x"274c0d3f", x"2fff254f", x"385a5b6f", x"f1260d3f", x"c8ce0000", x"f4880000", x"94a00000", x"ca5a8c20", x"c6be221a", x"73fd2787", x"c2e61309", x"929023e5"),
	(x"35a40000", x"8d0b0000", x"999d0000", x"c91e3440", x"c4403bb6", x"75b5c30c", x"db2fa3c7", x"70dbf437", x"2ee60000", x"b8c30000", x"3cf50000", x"198a8ec0", x"1edf12a2", x"eb5a975d", x"ea7315bd", x"45ca6b72"),
	(x"d38c0000", x"c1400000", x"31c80000", x"1ace36a0", x"1c210b0e", x"ed1273d6", x"f3baa573", x"a781bca0", x"de230000", x"e1e00000", x"79770000", x"f8078e00", x"25b21493", x"29b7c1c4", x"2193eba1", x"136ddaed"),
	(x"90a40000", x"bc5b0000", x"6d6e0000", x"0bdd4800", x"b728224a", x"ecc64a4f", x"759e1063", x"4cf701d1", x"36e70000", x"c9350000", x"d7980000", x"a32fa000", x"5a34515e", x"561c7179", x"310ab488", x"a074fe54"),
	(x"768c0000", x"f0100000", x"c53b0000", x"d80d4ae0", x"6f4912f2", x"7461fa95", x"5d0b16d7", x"9bad4946", x"c6220000", x"90160000", x"921a0000", x"42a2a0c0", x"6159576f", x"94f127e0", x"faea4a94", x"f6d34fcb"),
	(x"60610000", x"e5780000", x"28ec0000", x"ea5048c0", x"8c45247b", x"2e2b1cd6", x"be7eee7f", x"1a50b04e", x"200a0000", x"dc5d0000", x"3a4f0000", x"9172a220", x"b93867d7", x"0c56973a", x"d27f4c20", x"2189075c"),
	(x"86490000", x"a9330000", x"80b90000", x"39804a20", x"542414c3", x"b68cac0c", x"96ebe8cb", x"cd0af8d9", x"d0cf0000", x"857e0000", x"7fcd0000", x"70ffa2e0", x"825561e6", x"cebbc1a3", x"199fb23c", x"772eb6c3"),
	(x"24950000", x"cb680000", x"dc330000", x"740d4ce0", x"cf8a4372", x"3dd08912", x"a7c8c4ea", x"0298750f", x"d5e10000", x"74f40000", x"508b0000", x"1cdda060", x"748e5b44", x"dba94628", x"42cf1f8e", x"fba2eb6d"),
	(x"c2bd0000", x"87230000", x"74660000", x"a7dd4e00", x"17eb73ca", x"a57739c8", x"8f5dc25e", x"d5c23d98", x"25240000", x"2dd70000", x"15090000", x"fd50a0a0", x"4fe35d75", x"194410b1", x"892fe192", x"ad055af2"),
	(x"d4500000", x"924b0000", x"99b10000", x"95804c20", x"f4e74543", x"ff3ddf8b", x"6c283af6", x"543fc490", x"c30c0000", x"619c0000", x"bd5c0000", x"2e80a240", x"97826dcd", x"81e3a06b", x"a1bae726", x"7a5f1265"),
	(x"32780000", x"de000000", x"31e40000", x"46504ec0", x"2c8675fb", x"679a6f51", x"44bd3c42", x"83658c07", x"33c90000", x"38bf0000", x"f8de0000", x"cf0da280", x"acef6bfc", x"430ef6f2", x"6a5a193a", x"2cf8a3fa"),
	(x"73a20000", x"019a0000", x"ea7d0000", x"b42f4860", x"99922850", x"61737d1e", x"065bbb65", x"172114e8", x"61d00000", x"03c70000", x"e1d60000", x"630da480", x"0c2c3a7c", x"0abf8575", x"9099cb07", x"b5cd9fb3"),
	(x"958a0000", x"4dd10000", x"42280000", x"67ff4a80", x"41f318e8", x"f9d4cdc4", x"2ecebdd1", x"c07b5c7f", x"91150000", x"5ae40000", x"a4540000", x"8280a440", x"37413c4d", x"c852d3ec", x"5b79351b", x"e36a2e2c"),
	(x"83670000", x"58b90000", x"afff0000", x"55a248a0", x"a2ff2e61", x"a39e2b87", x"cdbb4579", x"4186a577", x"773d0000", x"16af0000", x"0c010000", x"5150a6a0", x"ef200cf5", x"50f56336", x"73ec33af", x"343066bb"),
	(x"654f0000", x"14f20000", x"07aa0000", x"86724a40", x"7a9e1ed9", x"3b399b5d", x"e52e43cd", x"96dcede0", x"87f80000", x"4f8c0000", x"49830000", x"b0dda660", x"d44d0ac4", x"921835af", x"b80ccdb3", x"6297d724"),
	(x"c7930000", x"76a90000", x"5b200000", x"cbff4c80", x"e1304968", x"b065be43", x"d40d6fec", x"594e6036", x"82d60000", x"be060000", x"66c50000", x"dcffa4e0", x"22963066", x"870ab224", x"e35c6001", x"ee1b8a8a"),
	(x"21bb0000", x"3ae20000", x"f3750000", x"182f4e60", x"395179d0", x"28c20e99", x"fc986958", x"8e1428a1", x"72130000", x"e7250000", x"23470000", x"3d72a420", x"19fb3657", x"45e7e4bd", x"28bc9e1d", x"b8bc3b15"),
	(x"37560000", x"2f8a0000", x"1ea20000", x"2a724c40", x"da5d4f59", x"7288e8da", x"1fed91f0", x"0fe9d1a9", x"943b0000", x"ab6e0000", x"8b120000", x"eea2a6c0", x"c19a06ef", x"dd405467", x"002998a9", x"6fe67382"),
	(x"d17e0000", x"63c10000", x"b6f70000", x"f9a24ea0", x"023c7fe1", x"ea2f5800", x"37789744", x"d8b3993e", x"64fe0000", x"f24d0000", x"ce900000", x"0f2fa600", x"faf700de", x"1fad02fe", x"cbc966b5", x"3941c21d"),
	(x"288b0000", x"0d770000", x"5db60000", x"1f991800", x"767042e8", x"dde1a2a3", x"5b06af40", x"19e93cbf", x"34150000", x"6bb40000", x"50a70000", x"4043d800", x"442925b1", x"51215aaf", x"f5c886bf", x"df46dbca"),
	(x"cea30000", x"413c0000", x"f5e30000", x"cc491ae0", x"ae117250", x"45461279", x"7393a9f4", x"ceb37428", x"c4d00000", x"32970000", x"15250000", x"a1ced8c0", x"7f442380", x"93cc0c36", x"3e2878a3", x"89e16a55"),
	(x"d84e0000", x"54540000", x"18340000", x"fe1418c0", x"4d1d44d9", x"1f0cf43a", x"90e6515c", x"4f4e8d20", x"22f80000", x"7edc0000", x"bd700000", x"721eda20", x"a7251338", x"0b6bbcec", x"16bd7e17", x"5ebb22c2"),
	(x"3e660000", x"181f0000", x"b0610000", x"2dc41a20", x"957c7461", x"87ab44e0", x"b87357e8", x"9814c5b7", x"d23d0000", x"27ff0000", x"f8f20000", x"9393dae0", x"9c481509", x"c986ea75", x"dd5d800b", x"081c935d"),
	(x"9cba0000", x"7a440000", x"eceb0000", x"60491ce0", x"0ed223d0", x"0cf761fe", x"89507bc9", x"57864861", x"d7130000", x"d6750000", x"d7b40000", x"ffb1d860", x"6a932fab", x"dc946dfe", x"860d2db9", x"8490cef3"),
	(x"7a920000", x"360f0000", x"44be0000", x"b3991e00", x"d6b31368", x"9450d124", x"a1c57d7d", x"80dc00f6", x"27d60000", x"8f560000", x"92360000", x"1e3cd8a0", x"51fe299a", x"1e793b67", x"4dedd3a5", x"d2377f6c"),
	(x"6c7f0000", x"23670000", x"a9690000", x"81c41c20", x"35bf25e1", x"ce1a3767", x"42b085d5", x"0121f9fe", x"c1fe0000", x"c31d0000", x"3a630000", x"cdecda40", x"899f1922", x"86de8bbd", x"6578d511", x"056d37fb"),
	(x"8a570000", x"6f2c0000", x"013c0000", x"52141ec0", x"edde1559", x"56bd87bd", x"6a258361", x"d67bb169", x"313b0000", x"9a3e0000", x"7fe10000", x"2c61da80", x"b2f21f13", x"4433dd24", x"ae982b0d", x"53ca8664"),
	(x"cb8d0000", x"b0b60000", x"daa50000", x"a06b1860", x"58ca48f2", x"505495f2", x"28c30446", x"423f2986", x"63220000", x"a1460000", x"66e90000", x"8061dc80", x"12314e93", x"0d82aea3", x"545bf930", x"caffba2d"),
	(x"2da50000", x"fcfd0000", x"72f00000", x"73bb1a80", x"80ab784a", x"c8f32528", x"005602f2", x"95656111", x"93e70000", x"f8650000", x"236b0000", x"61ecdc40", x"295c48a2", x"cf6ff83a", x"9fbb072c", x"9c580bb2"),
	(x"3b480000", x"e9950000", x"9f270000", x"41e618a0", x"63a74ec3", x"92b9c36b", x"e323fa5a", x"14989819", x"75cf0000", x"b42e0000", x"8b3e0000", x"b23cdea0", x"f13d781a", x"57c848e0", x"b72e0198", x"4b024325"),
	(x"dd600000", x"a5de0000", x"37720000", x"92361a40", x"bbc67e7b", x"0a1e73b1", x"cbb6fcee", x"c3c2d08e", x"850a0000", x"ed0d0000", x"cebc0000", x"53b1de60", x"ca507e2b", x"95251e79", x"7cceff84", x"1da5f2ba"),
	(x"7fbc0000", x"c7850000", x"6bf80000", x"dfbb1c80", x"206829ca", x"814256af", x"fa95d0cf", x"0c505d58", x"80240000", x"1c870000", x"e1fa0000", x"3f93dce0", x"3c8b4489", x"803799f2", x"279e5236", x"9129af14"),
	(x"99940000", x"8bce0000", x"c3ad0000", x"0c6b1e60", x"f8091972", x"19e5e675", x"d200d67b", x"db0a15cf", x"70e10000", x"45a40000", x"a4780000", x"de1edc20", x"07e642b8", x"42dacf6b", x"ec7eac2a", x"c78e1e8b"),
	(x"8f790000", x"9ea60000", x"2e7a0000", x"3e361c40", x"1b052ffb", x"43af0036", x"31752ed3", x"5af7ecc7", x"96c90000", x"09ef0000", x"0c2d0000", x"0dcedec0", x"df877200", x"da7d7fb1", x"c4ebaa9e", x"10d4561c"),
	(x"69510000", x"d2ed0000", x"862f0000", x"ede61ea0", x"c3641f43", x"db08b0ec", x"19e02867", x"8dada450", x"660c0000", x"50cc0000", x"49af0000", x"ec43de00", x"e4ea7431", x"18902928", x"0f0b5482", x"4673e783"),
	(x"2a790000", x"aff60000", x"da890000", x"fcf56000", x"686d3607", x"dadc8975", x"9fc49d77", x"66db1921", x"8ec80000", x"78190000", x"e7400000", x"b76bf000", x"9b6c31fc", x"673b9995", x"1f920bab", x"f56ac33a"),
	(x"cc510000", x"e3bd0000", x"72dc0000", x"2f2562e0", x"b00c06bf", x"427b39af", x"b7519bc3", x"b18151b6", x"7e0d0000", x"213a0000", x"a2c20000", x"56e6f0c0", x"a00137cd", x"a5d6cf0c", x"d472f5b7", x"a3cd72a5"),
	(x"dabc0000", x"f6d50000", x"9f0b0000", x"1d7860c0", x"53003036", x"1831dfec", x"5424636b", x"307ca8be", x"98250000", x"6d710000", x"0a970000", x"8536f220", x"78600775", x"3d717fd6", x"fce7f303", x"74973a32"),
	(x"3c940000", x"ba9e0000", x"375e0000", x"cea86220", x"8b61008e", x"80966f36", x"7cb165df", x"e726e029", x"68e00000", x"34520000", x"4f150000", x"64bbf2e0", x"430d0144", x"ff9c294f", x"37070d1f", x"22308bad"),
	(x"9e480000", x"d8c50000", x"6bd40000", x"832564e0", x"10cf573f", x"0bca4a28", x"4d9249fe", x"28b46dff", x"6dce0000", x"c5d80000", x"60530000", x"0899f060", x"b5d63be6", x"ea8eaec4", x"6c57a0ad", x"aebcd603"),
	(x"78600000", x"948e0000", x"c3810000", x"50f56600", x"c8ae6787", x"936dfaf2", x"65074f4a", x"ffee2568", x"9d0b0000", x"9cfb0000", x"25d10000", x"e914f0a0", x"8ebb3dd7", x"2863f85d", x"a7b75eb1", x"f81b679c"),
	(x"6e8d0000", x"81e60000", x"2e560000", x"62a86420", x"2ba2510e", x"c9271cb1", x"8672b7e2", x"7e13dc60", x"7b230000", x"d0b00000", x"8d840000", x"3ac4f240", x"56da0d6f", x"b0c44887", x"8f225805", x"2f412f0b"),
	(x"88a50000", x"cdad0000", x"86030000", x"b17866c0", x"f3c361b6", x"5180ac6b", x"aee7b156", x"a94994f7", x"8be60000", x"89930000", x"c8060000", x"db49f280", x"6db70b5e", x"72291e1e", x"44c2a619", x"79e69e94"),
	(x"c97f0000", x"12370000", x"5d9a0000", x"43076060", x"46d73c1d", x"5769be24", x"ec013671", x"3d0d0c18", x"d9ff0000", x"b2eb0000", x"d10e0000", x"7749f480", x"cd745ade", x"3b986d99", x"be017424", x"e0d3a2dd"),
	(x"2f570000", x"5e7c0000", x"f5cf0000", x"90d76280", x"9eb60ca5", x"cfce0efe", x"c49430c5", x"ea57448f", x"293a0000", x"ebc80000", x"948c0000", x"96c4f440", x"f6195cef", x"f9753b00", x"75e18a38", x"b6741342"),
	(x"39ba0000", x"4b140000", x"18180000", x"a28a60a0", x"7dba3a2c", x"9584e8bd", x"27e1c86d", x"6baabd87", x"cf120000", x"a7830000", x"3cd90000", x"4514f6a0", x"2e786c57", x"61d28bda", x"5d748c8c", x"612e5bd5"),
	(x"df920000", x"075f0000", x"b04d0000", x"715a6240", x"a5db0a94", x"0d235867", x"0f74ced9", x"bcf0f510", x"3fd70000", x"fea00000", x"795b0000", x"a499f660", x"15156a66", x"a33fdd43", x"96947290", x"3789ea4a"),
	(x"7d4e0000", x"65040000", x"ecc70000", x"3cd76480", x"3e755d25", x"867f7d79", x"3e57e2f8", x"736278c6", x"3af90000", x"0f2a0000", x"561d0000", x"c8bbf4e0", x"e3ce50c4", x"b62d5ac8", x"cdc4df22", x"bb05b7e4"),
	(x"9b660000", x"294f0000", x"44920000", x"ef076660", x"e6146d9d", x"1ed8cda3", x"16c2e44c", x"a4383051", x"ca3c0000", x"56090000", x"139f0000", x"2936f420", x"d8a356f5", x"74c00c51", x"0624213e", x"eda2067b"),
	(x"8d8b0000", x"3c270000", x"a9450000", x"dd5a6440", x"05185b14", x"44922be0", x"f5b71ce4", x"25c5c959", x"2c140000", x"1a420000", x"bbca0000", x"fae6f6c0", x"00c2664d", x"ec67bc8b", x"2eb1278a", x"3af84eec"),
	(x"6ba30000", x"706c0000", x"01100000", x"0e8a66a0", x"dd796bac", x"dc359b3a", x"dd221a50", x"f29f81ce", x"dcd10000", x"43610000", x"fe480000", x"1b6bf600", x"3baf607c", x"2e8aea12", x"e551d996", x"6c5fff73"),
	(x"8c3a0000", x"da980000", x"607f0000", x"54078800", x"85714513", x"6006b243", x"db50399c", x"8a58e6a4", x"1e6c0000", x"c4420000", x"8a2e0000", x"bcb6b800", x"2c4413b6", x"8bfdd3da", x"6a0c1bc8", x"b99dc2eb"),
	(x"6a120000", x"96d30000", x"c82a0000", x"87d78ae0", x"5d1075ab", x"f8a10299", x"f3c53f28", x"5d02ae33", x"eea90000", x"9d610000", x"cfac0000", x"5d3bb8c0", x"17291587", x"49108543", x"a1ece5d4", x"ef3a7374"),
	(x"7cff0000", x"83bb0000", x"25fd0000", x"b58a88c0", x"be1c4322", x"a2ebe4da", x"10b0c780", x"dcff573b", x"08810000", x"d12a0000", x"67f90000", x"8eebba20", x"cf48253f", x"d1b73599", x"8979e360", x"38603be3"),
	(x"9ad70000", x"cff00000", x"8da80000", x"665a8a20", x"667d739a", x"3a4c5400", x"3825c134", x"0ba51fac", x"f8440000", x"88090000", x"227b0000", x"6f66bae0", x"f425230e", x"135a6300", x"42991d7c", x"6ec78a7c"),
	(x"380b0000", x"adab0000", x"d1220000", x"2bd78ce0", x"fdd3242b", x"b110711e", x"0906ed15", x"c437927a", x"fd6a0000", x"79830000", x"0d3d0000", x"0344b860", x"02fe19ac", x"0648e48b", x"19c9b0ce", x"e24bd7d2"),
	(x"de230000", x"e1e00000", x"79770000", x"f8078e00", x"25b21493", x"29b7c1c4", x"2193eba1", x"136ddaed", x"0daf0000", x"20a00000", x"48bf0000", x"e2c9b8a0", x"39931f9d", x"c4a5b212", x"d2294ed2", x"b4ec664d"),
	(x"c8ce0000", x"f4880000", x"94a00000", x"ca5a8c20", x"c6be221a", x"73fd2787", x"c2e61309", x"929023e5", x"eb870000", x"6ceb0000", x"e0ea0000", x"3119ba40", x"e1f22f25", x"5c0202c8", x"fabc4866", x"63b62eda"),
	(x"2ee60000", x"b8c30000", x"3cf50000", x"198a8ec0", x"1edf12a2", x"eb5a975d", x"ea7315bd", x"45ca6b72", x"1b420000", x"35c80000", x"a5680000", x"d094ba80", x"da9f2914", x"9eef5451", x"315cb67a", x"35119f45"),
	(x"6f3c0000", x"67590000", x"e76c0000", x"ebf58860", x"abcb4f09", x"edb38512", x"a895929a", x"d18ef39d", x"495b0000", x"0eb00000", x"bc600000", x"7c94bc80", x"7a5c7894", x"d75e27d6", x"cb9f6447", x"ac24a30c"),
	(x"89140000", x"2b120000", x"4f390000", x"38258a80", x"73aa7fb1", x"751435c8", x"8000942e", x"06d4bb0a", x"b99e0000", x"57930000", x"f9e20000", x"9d19bc40", x"41317ea5", x"15b3714f", x"007f9a5b", x"fa831293"),
	(x"9ff90000", x"3e7a0000", x"a2ee0000", x"0a7888a0", x"90a64938", x"2f5ed38b", x"63756c86", x"87294202", x"5fb60000", x"1bd80000", x"51b70000", x"4ec9bea0", x"99504e1d", x"8d14c195", x"28ea9cef", x"2dd95a04"),
	(x"79d10000", x"72310000", x"0abb0000", x"d9a88a40", x"48c77980", x"b7f96351", x"4be06a32", x"50730a95", x"af730000", x"42fb0000", x"14350000", x"af44be60", x"a23d482c", x"4ff9970c", x"e30a62f3", x"7b7eeb9b"),
	(x"db0d0000", x"106a0000", x"56310000", x"94258c80", x"d3692e31", x"3ca5464f", x"7ac34613", x"9fe18743", x"aa5d0000", x"b3710000", x"3b730000", x"c366bce0", x"54e6728e", x"5aeb1087", x"b85acf41", x"f7f2b635"),
	(x"3d250000", x"5c210000", x"fe640000", x"47f58e60", x"0b081e89", x"a402f695", x"525640a7", x"48bbcfd4", x"5a980000", x"ea520000", x"7ef10000", x"22ebbc20", x"6f8b74bf", x"9806461e", x"73ba315d", x"a15507aa"),
	(x"2bc80000", x"49490000", x"13b30000", x"75a88c40", x"e8042800", x"fe4810d6", x"b123b80f", x"c94636dc", x"bcb00000", x"a6190000", x"d6a40000", x"f13bbec0", x"b7ea4407", x"00a1f6c4", x"5b2f37e9", x"760f4f3d"),
	(x"cde00000", x"05020000", x"bbe60000", x"a6788ea0", x"306518b8", x"66efa00c", x"99b6bebb", x"1e1c7e4b", x"4c750000", x"ff3a0000", x"93260000", x"10b6be00", x"8c874236", x"c24ca05d", x"90cfc9f5", x"20a8fea2"),
	(x"8ec80000", x"78190000", x"e7400000", x"b76bf000", x"9b6c31fc", x"673b9995", x"1f920bab", x"f56ac33a", x"a4b10000", x"d7ef0000", x"3dc90000", x"4b9e9000", x"f30107fb", x"bde710e0", x"805696dc", x"93b1da1b"),
	(x"68e00000", x"34520000", x"4f150000", x"64bbf2e0", x"430d0144", x"ff9c294f", x"37070d1f", x"22308bad", x"54740000", x"8ecc0000", x"784b0000", x"aa1390c0", x"c86c01ca", x"7f0a4679", x"4bb668c0", x"c5166b84"),
	(x"7e0d0000", x"213a0000", x"a2c20000", x"56e6f0c0", x"a00137cd", x"a5d6cf0c", x"d472f5b7", x"a3cd72a5", x"b25c0000", x"c2870000", x"d01e0000", x"79c39220", x"100d3172", x"e7adf6a3", x"63236e74", x"124c2313"),
	(x"98250000", x"6d710000", x"0a970000", x"8536f220", x"78600775", x"3d717fd6", x"fce7f303", x"74973a32", x"42990000", x"9ba40000", x"959c0000", x"984e92e0", x"2b603743", x"2540a03a", x"a8c39068", x"44eb928c"),
	(x"3af90000", x"0f2a0000", x"561d0000", x"c8bbf4e0", x"e3ce50c4", x"b62d5ac8", x"cdc4df22", x"bb05b7e4", x"47b70000", x"6a2e0000", x"bada0000", x"f46c9060", x"ddbb0de1", x"305227b1", x"f3933dda", x"c867cf22"),
	(x"dcd10000", x"43610000", x"fe480000", x"1b6bf600", x"3baf607c", x"2e8aea12", x"e551d996", x"6c5fff73", x"b7720000", x"330d0000", x"ff580000", x"15e190a0", x"e6d60bd0", x"f2bf7128", x"3873c3c6", x"9ec07ebd"),
	(x"ca3c0000", x"56090000", x"139f0000", x"2936f420", x"d8a356f5", x"74c00c51", x"0624213e", x"eda2067b", x"515a0000", x"7f460000", x"570d0000", x"c6319240", x"3eb73b68", x"6a18c1f2", x"10e6c572", x"499a362a"),
	(x"2c140000", x"1a420000", x"bbca0000", x"fae6f6c0", x"00c2664d", x"ec67bc8b", x"2eb1278a", x"3af84eec", x"a19f0000", x"26650000", x"128f0000", x"27bc9280", x"05da3d59", x"a8f5976b", x"db063b6e", x"1f3d87b5"),
	(x"6dce0000", x"c5d80000", x"60530000", x"0899f060", x"b5d63be6", x"ea8eaec4", x"6c57a0ad", x"aebcd603", x"f3860000", x"1d1d0000", x"0b870000", x"8bbc9480", x"a5196cd9", x"e144e4ec", x"21c5e953", x"8608bbfc"),
	(x"8be60000", x"89930000", x"c8060000", x"db49f280", x"6db70b5e", x"72291e1e", x"44c2a619", x"79e69e94", x"03430000", x"443e0000", x"4e050000", x"6a319440", x"9e746ae8", x"23a9b275", x"ea25174f", x"d0af0a63"),
	(x"9d0b0000", x"9cfb0000", x"25d10000", x"e914f0a0", x"8ebb3dd7", x"2863f85d", x"a7b75eb1", x"f81b679c", x"e56b0000", x"08750000", x"e6500000", x"b9e196a0", x"46155a50", x"bb0e02af", x"c2b011fb", x"07f542f4"),
	(x"7b230000", x"d0b00000", x"8d840000", x"3ac4f240", x"56da0d6f", x"b0c44887", x"8f225805", x"2f412f0b", x"15ae0000", x"51560000", x"a3d20000", x"586c9660", x"7d785c61", x"79e35436", x"0950efe7", x"5152f36b"),
	(x"d9ff0000", x"b2eb0000", x"d10e0000", x"7749f480", x"cd745ade", x"3b986d99", x"be017424", x"e0d3a2dd", x"10800000", x"a0dc0000", x"8c940000", x"344e94e0", x"8ba366c3", x"6cf1d3bd", x"52004255", x"dddeaec5"),
	(x"3fd70000", x"fea00000", x"795b0000", x"a499f660", x"15156a66", x"a33fdd43", x"96947290", x"3789ea4a", x"e0450000", x"f9ff0000", x"c9160000", x"d5c39420", x"b0ce60f2", x"ae1c8524", x"99e0bc49", x"8b791f5a"),
	(x"293a0000", x"ebc80000", x"948c0000", x"96c4f440", x"f6195cef", x"f9753b00", x"75e18a38", x"b6741342", x"066d0000", x"b5b40000", x"61430000", x"061396c0", x"68af504a", x"36bb35fe", x"b175bafd", x"5c2357cd"),
	(x"cf120000", x"a7830000", x"3cd90000", x"4514f6a0", x"2e786c57", x"61d28bda", x"5d748c8c", x"612e5bd5", x"f6a80000", x"ec970000", x"24c10000", x"e79e9600", x"53c2567b", x"f4566367", x"7a9544e1", x"0a84e652"),
	(x"36e70000", x"c9350000", x"d7980000", x"a32fa000", x"5a34515e", x"561c7179", x"310ab488", x"a074fe54", x"a6430000", x"756e0000", x"baf60000", x"a8f2e800", x"ed1c7314", x"bada3b36", x"4494a4eb", x"ec83ff85"),
	(x"d0cf0000", x"857e0000", x"7fcd0000", x"70ffa2e0", x"825561e6", x"cebbc1a3", x"199fb23c", x"772eb6c3", x"56860000", x"2c4d0000", x"ff740000", x"497fe8c0", x"d6717525", x"78376daf", x"8f745af7", x"ba244e1a"),
	(x"c6220000", x"90160000", x"921a0000", x"42a2a0c0", x"6159576f", x"94f127e0", x"faea4a94", x"f6d34fcb", x"b0ae0000", x"60060000", x"57210000", x"9aafea20", x"0e10459d", x"e090dd75", x"a7e15c43", x"6d7e068d"),
	(x"200a0000", x"dc5d0000", x"3a4f0000", x"9172a220", x"b93867d7", x"0c56973a", x"d27f4c20", x"2189075c", x"406b0000", x"39250000", x"12a30000", x"7b22eae0", x"357d43ac", x"227d8bec", x"6c01a25f", x"3bd9b712"),
	(x"82d60000", x"be060000", x"66c50000", x"dcffa4e0", x"22963066", x"870ab224", x"e35c6001", x"ee1b8a8a", x"45450000", x"c8af0000", x"3de50000", x"1700e860", x"c3a6790e", x"376f0c67", x"37510fed", x"b755eabc"),
	(x"64fe0000", x"f24d0000", x"ce900000", x"0f2fa600", x"faf700de", x"1fad02fe", x"cbc966b5", x"3941c21d", x"b5800000", x"918c0000", x"78670000", x"f68de8a0", x"f8cb7f3f", x"f5825afe", x"fcb1f1f1", x"e1f25b23"),
	(x"72130000", x"e7250000", x"23470000", x"3d72a420", x"19fb3657", x"45e7e4bd", x"28bc9e1d", x"b8bc3b15", x"53a80000", x"ddc70000", x"d0320000", x"255dea40", x"20aa4f87", x"6d25ea24", x"d424f745", x"36a813b4"),
	(x"943b0000", x"ab6e0000", x"8b120000", x"eea2a6c0", x"c19a06ef", x"dd405467", x"002998a9", x"6fe67382", x"a36d0000", x"84e40000", x"95b00000", x"c4d0ea80", x"1bc749b6", x"afc8bcbd", x"1fc40959", x"600fa22b"),
	(x"d5e10000", x"74f40000", x"508b0000", x"1cdda060", x"748e5b44", x"dba94628", x"42cf1f8e", x"fba2eb6d", x"f1740000", x"bf9c0000", x"8cb80000", x"68d0ec80", x"bb041836", x"e679cf3a", x"e507db64", x"f93a9e62"),
	(x"33c90000", x"38bf0000", x"f8de0000", x"cf0da280", x"acef6bfc", x"430ef6f2", x"6a5a193a", x"2cf8a3fa", x"01b10000", x"e6bf0000", x"c93a0000", x"895dec40", x"80691e07", x"249499a3", x"2ee72578", x"af9d2ffd"),
	(x"25240000", x"2dd70000", x"15090000", x"fd50a0a0", x"4fe35d75", x"194410b1", x"892fe192", x"ad055af2", x"e7990000", x"aaf40000", x"616f0000", x"5a8deea0", x"58082ebf", x"bc332979", x"067223cc", x"78c7676a"),
	(x"c30c0000", x"619c0000", x"bd5c0000", x"2e80a240", x"97826dcd", x"81e3a06b", x"a1bae726", x"7a5f1265", x"175c0000", x"f3d70000", x"24ed0000", x"bb00ee60", x"6365288e", x"7ede7fe0", x"cd92ddd0", x"2e60d6f5"),
	(x"61d00000", x"03c70000", x"e1d60000", x"630da480", x"0c2c3a7c", x"0abf8575", x"9099cb07", x"b5cd9fb3", x"12720000", x"025d0000", x"0bab0000", x"d722ece0", x"95be122c", x"6bccf86b", x"96c27062", x"a2ec8b5b"),
	(x"87f80000", x"4f8c0000", x"49830000", x"b0dda660", x"d44d0ac4", x"921835af", x"b80ccdb3", x"6297d724", x"e2b70000", x"5b7e0000", x"4e290000", x"36afec20", x"aed3141d", x"a921aef2", x"5d228e7e", x"f44b3ac4"),
	(x"91150000", x"5ae40000", x"a4540000", x"8280a440", x"37413c4d", x"c852d3ec", x"5b79351b", x"e36a2e2c", x"049f0000", x"17350000", x"e67c0000", x"e57feec0", x"76b224a5", x"31861e28", x"75b788ca", x"23117253"),
	(x"773d0000", x"16af0000", x"0c010000", x"5150a6a0", x"ef200cf5", x"50f56336", x"73ec33af", x"343066bb", x"f45a0000", x"4e160000", x"a3fe0000", x"04f2ee00", x"4ddf2294", x"f36b48b1", x"be5776d6", x"75b6c3cc"),
	(x"34150000", x"6bb40000", x"50a70000", x"4043d800", x"442925b1", x"51215aaf", x"f5c886bf", x"df46dbca", x"1c9e0000", x"66c30000", x"0d110000", x"5fdac000", x"32596759", x"8cc0f80c", x"aece29ff", x"c6afe775"),
	(x"d23d0000", x"27ff0000", x"f8f20000", x"9393dae0", x"9c481509", x"c986ea75", x"dd5d800b", x"081c935d", x"ec5b0000", x"3fe00000", x"48930000", x"be57c0c0", x"09346168", x"4e2dae95", x"652ed7e3", x"900856ea"),
	(x"c4d00000", x"32970000", x"15250000", x"a1ced8c0", x"7f442380", x"93cc0c36", x"3e2878a3", x"89e16a55", x"0a730000", x"73ab0000", x"e0c60000", x"6d87c220", x"d15551d0", x"d68a1e4f", x"4dbbd157", x"47521e7d"),
	(x"22f80000", x"7edc0000", x"bd700000", x"721eda20", x"a7251338", x"0b6bbcec", x"16bd7e17", x"5ebb22c2", x"fab60000", x"2a880000", x"a5440000", x"8c0ac2e0", x"ea3857e1", x"146748d6", x"865b2f4b", x"11f5afe2"),
	(x"80240000", x"1c870000", x"e1fa0000", x"3f93dce0", x"3c8b4489", x"803799f2", x"279e5236", x"9129af14", x"ff980000", x"db020000", x"8a020000", x"e028c060", x"1ce36d43", x"0175cf5d", x"dd0b82f9", x"9d79f24c"),
	(x"660c0000", x"50cc0000", x"49af0000", x"ec43de00", x"e4ea7431", x"18902928", x"0f0b5482", x"4673e783", x"0f5d0000", x"82210000", x"cf800000", x"01a5c0a0", x"278e6b72", x"c39899c4", x"16eb7ce5", x"cbde43d3"),
	(x"70e10000", x"45a40000", x"a4780000", x"de1edc20", x"07e642b8", x"42dacf6b", x"ec7eac2a", x"c78e1e8b", x"e9750000", x"ce6a0000", x"67d50000", x"d275c240", x"ffef5bca", x"5b3f291e", x"3e7e7a51", x"1c840b44"),
	(x"96c90000", x"09ef0000", x"0c2d0000", x"0dcedec0", x"df877200", x"da7d7fb1", x"c4ebaa9e", x"10d4561c", x"19b00000", x"97490000", x"22570000", x"33f8c280", x"c4825dfb", x"99d27f87", x"f59e844d", x"4a23badb"),
	(x"d7130000", x"d6750000", x"d7b40000", x"ffb1d860", x"6a932fab", x"dc946dfe", x"860d2db9", x"8490cef3", x"4ba90000", x"ac310000", x"3b5f0000", x"9ff8c480", x"64410c7b", x"d0630c00", x"0f5d5670", x"d3168692"),
	(x"313b0000", x"9a3e0000", x"7fe10000", x"2c61da80", x"b2f21f13", x"4433dd24", x"ae982b0d", x"53ca8664", x"bb6c0000", x"f5120000", x"7edd0000", x"7e75c440", x"5f2c0a4a", x"128e5a99", x"c4bda86c", x"85b1370d"),
	(x"27d60000", x"8f560000", x"92360000", x"1e3cd8a0", x"51fe299a", x"1e793b67", x"4dedd3a5", x"d2377f6c", x"5d440000", x"b9590000", x"d6880000", x"ada5c6a0", x"874d3af2", x"8a29ea43", x"ec28aed8", x"52eb7f9a"),
	(x"c1fe0000", x"c31d0000", x"3a630000", x"cdecda40", x"899f1922", x"86de8bbd", x"6578d511", x"056d37fb", x"ad810000", x"e07a0000", x"930a0000", x"4c28c660", x"bc203cc3", x"48c4bcda", x"27c850c4", x"044cce05"),
	(x"63220000", x"a1460000", x"66e90000", x"8061dc80", x"12314e93", x"0d82aea3", x"545bf930", x"caffba2d", x"a8af0000", x"11f00000", x"bc4c0000", x"200ac4e0", x"4afb0661", x"5dd63b51", x"7c98fd76", x"88c093ab"),
	(x"850a0000", x"ed0d0000", x"cebc0000", x"53b1de60", x"ca507e2b", x"95251e79", x"7cceff84", x"1da5f2ba", x"586a0000", x"48d30000", x"f9ce0000", x"c187c420", x"71960050", x"9f3b6dc8", x"b778036a", x"de672234"),
	(x"93e70000", x"f8650000", x"236b0000", x"61ecdc40", x"295c48a2", x"cf6ff83a", x"9fbb072c", x"9c580bb2", x"be420000", x"04980000", x"519b0000", x"1257c6c0", x"a9f730e8", x"079cdd12", x"9fed05de", x"093d6aa3"),
	(x"75cf0000", x"b42e0000", x"8b3e0000", x"b23cdea0", x"f13d781a", x"57c848e0", x"b72e0198", x"4b024325", x"4e870000", x"5dbb0000", x"14190000", x"f3dac600", x"929a36d9", x"c5718b8b", x"540dfbc2", x"5f9adb3c")
    ),(
	(x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000"),
	(x"033d0000", x"08b30000", x"f33a0000", x"3ac20007", x"51298a50", x"6b6e661f", x"0ea5cfe3", x"e6da7ffe", x"a8da0000", x"96be0000", x"5c1d0000", x"07da0002", x"7d669583", x"1f98708a", x"bb668808", x"da878000"),
	(x"a8da0000", x"96be0000", x"5c1d0000", x"07da0002", x"7d669583", x"1f98708a", x"bb668808", x"da878000", x"abe70000", x"9e0d0000", x"af270000", x"3d180005", x"2c4f1fd3", x"74f61695", x"b5c347eb", x"3c5dfffe"),
	(x"abe70000", x"9e0d0000", x"af270000", x"3d180005", x"2c4f1fd3", x"74f61695", x"b5c347eb", x"3c5dfffe", x"033d0000", x"08b30000", x"f33a0000", x"3ac20007", x"51298a50", x"6b6e661f", x"0ea5cfe3", x"e6da7ffe"),
	(x"01930000", x"e7820000", x"edfb0000", x"cf0c000b", x"8dd08d58", x"bca3b42e", x"063661e1", x"536f9e7b", x"92280000", x"dc850000", x"57fa0000", x"56dc0003", x"bae92316", x"5aefa30c", x"90cef752", x"7b1675d7"),
	(x"02ae0000", x"ef310000", x"1ec10000", x"f5ce000c", x"dcf90708", x"d7cdd231", x"0893ae02", x"b5b5e185", x"3af20000", x"4a3b0000", x"0be70000", x"51060001", x"c78fb695", x"4577d386", x"2ba87f5a", x"a191f5d7"),
	(x"a9490000", x"713c0000", x"b1e60000", x"c8d60009", x"f0b618db", x"a33bc4a4", x"bd50e9e9", x"89e81e7b", x"39cf0000", x"42880000", x"f8dd0000", x"6bc40006", x"96a63cc5", x"2e19b599", x"250db0b9", x"474b8a29"),
	(x"aa740000", x"798f0000", x"42dc0000", x"f214000e", x"a19f928b", x"c855a2bb", x"b3f5260a", x"6f326185", x"91150000", x"d4360000", x"a4c00000", x"6c1e0004", x"ebc0a946", x"3181c513", x"9e6b38b1", x"9dcc0a29"),
	(x"92280000", x"dc850000", x"57fa0000", x"56dc0003", x"bae92316", x"5aefa30c", x"90cef752", x"7b1675d7", x"93bb0000", x"3b070000", x"ba010000", x"99d00008", x"3739ae4e", x"e64c1722", x"96f896b3", x"2879ebac"),
	(x"91150000", x"d4360000", x"a4c00000", x"6c1e0004", x"ebc0a946", x"3181c513", x"9e6b38b1", x"9dcc0a29", x"3b610000", x"adb90000", x"e61c0000", x"9e0a000a", x"4a5f3bcd", x"f9d467a8", x"2d9e1ebb", x"f2fe6bac"),
	(x"3af20000", x"4a3b0000", x"0be70000", x"51060001", x"c78fb695", x"4577d386", x"2ba87f5a", x"a191f5d7", x"385c0000", x"a50a0000", x"15260000", x"a4c8000d", x"1b76b19d", x"92ba01b7", x"233bd158", x"14241452"),
	(x"39cf0000", x"42880000", x"f8dd0000", x"6bc40006", x"96a63cc5", x"2e19b599", x"250db0b9", x"474b8a29", x"90860000", x"33b40000", x"493b0000", x"a312000f", x"6610241e", x"8d22713d", x"985d5950", x"cea39452"),
	(x"93bb0000", x"3b070000", x"ba010000", x"99d00008", x"3739ae4e", x"e64c1722", x"96f896b3", x"2879ebac", x"01930000", x"e7820000", x"edfb0000", x"cf0c000b", x"8dd08d58", x"bca3b42e", x"063661e1", x"536f9e7b"),
	(x"90860000", x"33b40000", x"493b0000", x"a312000f", x"6610241e", x"8d22713d", x"985d5950", x"cea39452", x"a9490000", x"713c0000", x"b1e60000", x"c8d60009", x"f0b618db", x"a33bc4a4", x"bd50e9e9", x"89e81e7b"),
	(x"3b610000", x"adb90000", x"e61c0000", x"9e0a000a", x"4a5f3bcd", x"f9d467a8", x"2d9e1ebb", x"f2fe6bac", x"aa740000", x"798f0000", x"42dc0000", x"f214000e", x"a19f928b", x"c855a2bb", x"b3f5260a", x"6f326185"),
	(x"385c0000", x"a50a0000", x"15260000", x"a4c8000d", x"1b76b19d", x"92ba01b7", x"233bd158", x"14241452", x"02ae0000", x"ef310000", x"1ec10000", x"f5ce000c", x"dcf90708", x"d7cdd231", x"0893ae02", x"b5b5e185"),
	(x"5fa80000", x"56030000", x"43ae0000", x"64f30013", x"257e86bf", x"1311944e", x"541e95bf", x"8ea4db69", x"00440000", x"7f480000", x"da7c0000", x"2a230001", x"3badc9cc", x"a9b69c87", x"030a9e60", x"be0a679e"),
	(x"5c950000", x"5eb00000", x"b0940000", x"5e310014", x"74570cef", x"787ff251", x"5abb5a5c", x"687ea497", x"a89e0000", x"e9f60000", x"86610000", x"2df90003", x"46cb5c4f", x"b62eec0d", x"b86c1668", x"648de79e"),
	(x"f7720000", x"c0bd0000", x"1fb30000", x"63290011", x"5818133c", x"0c89e4c4", x"ef781db7", x"54235b69", x"aba30000", x"e1450000", x"755b0000", x"173b0004", x"17e2d61f", x"dd408a12", x"b6c9d98b", x"82579860"),
	(x"f44f0000", x"c80e0000", x"ec890000", x"59eb0016", x"0931996c", x"67e782db", x"e1ddd254", x"b2f92497", x"03790000", x"77fb0000", x"29460000", x"10e10006", x"6a84439c", x"c2d8fa98", x"0daf5183", x"58d01860"),
	(x"5e3b0000", x"b1810000", x"ae550000", x"abff0018", x"a8ae0be7", x"afb22060", x"5228f45e", x"ddcb4512", x"926c0000", x"a3cd0000", x"8d860000", x"7cff0002", x"8144eada", x"f3593f8b", x"93c46932", x"c51c1249"),
	(x"5d060000", x"b9320000", x"5d6f0000", x"913d001f", x"f98781b7", x"c4dc467f", x"5c8d3bbd", x"3b113aec", x"3ab60000", x"35730000", x"d19b0000", x"7b250000", x"fc227f59", x"ecc14f01", x"28a2e13a", x"1f9b9249"),
	(x"f6e10000", x"273f0000", x"f2480000", x"ac25001a", x"d5c89e64", x"b02a50ea", x"e94e7c56", x"074cc512", x"398b0000", x"3dc00000", x"22a10000", x"41e70007", x"ad0bf509", x"87af291e", x"26072ed9", x"f941edb7"),
	(x"f5dc0000", x"2f8c0000", x"01720000", x"96e7001d", x"84e11434", x"db4436f5", x"e7ebb3b5", x"e196baec", x"91510000", x"ab7e0000", x"7ebc0000", x"463d0005", x"d06d608a", x"98375994", x"9d61a6d1", x"23c66db7"),
	(x"cd800000", x"8a860000", x"14540000", x"322f0010", x"9f97a5a9", x"49fe3742", x"c4d062ed", x"f5b2aebe", x"93ff0000", x"444f0000", x"607d0000", x"b3f30009", x"0c946782", x"4ffa8ba5", x"95f208d3", x"96738c32"),
	(x"cebd0000", x"82350000", x"e76e0000", x"08ed0017", x"cebe2ff9", x"2290515d", x"ca75ad0e", x"1368d140", x"3b250000", x"d2f10000", x"3c600000", x"b429000b", x"71f2f201", x"5062fb2f", x"2e9480db", x"4cf40c32"),
	(x"655a0000", x"1c380000", x"48490000", x"35f50012", x"e2f1302a", x"566647c8", x"7fb6eae5", x"2f352ebe", x"38180000", x"da420000", x"cf5a0000", x"8eeb000c", x"20db7851", x"3b0c9d30", x"20314f38", x"aa2e73cc"),
	(x"66670000", x"148b0000", x"bb730000", x"0f370015", x"b3d8ba7a", x"3d0821d7", x"71132506", x"c9ef5140", x"90c20000", x"4cfc0000", x"93470000", x"8931000e", x"5dbdedd2", x"2494edba", x"9b57c730", x"70a9f3cc"),
	(x"cc130000", x"6d040000", x"f9af0000", x"fd23001b", x"124728f1", x"f55d836c", x"c2e6030c", x"a6dd30c5", x"01d70000", x"98ca0000", x"37870000", x"e52f000a", x"b67d4494", x"151528a9", x"053cff81", x"ed65f9e5"),
	(x"cf2e0000", x"65b70000", x"0a950000", x"c7e1001c", x"436ea2a1", x"9e33e573", x"cc43ccef", x"40074f3b", x"a90d0000", x"0e740000", x"6b9a0000", x"e2f50008", x"cb1bd117", x"0a8d5823", x"be5a7789", x"37e279e5"),
	(x"64c90000", x"fbba0000", x"a5b20000", x"faf90019", x"6f21bd72", x"eac5f3e6", x"79808b04", x"7c5ab0c5", x"aa300000", x"06c70000", x"98a00000", x"d837000f", x"9a325b47", x"61e33e3c", x"b0ffb86a", x"d138061b"),
	(x"67f40000", x"f3090000", x"56880000", x"c03b001e", x"3e083722", x"81ab95f9", x"772544e7", x"9a80cf3b", x"02ea0000", x"90790000", x"c4bd0000", x"dfed000d", x"e754cec4", x"7e7b4eb6", x"0b993062", x"0bbf861b"),
	(x"00440000", x"7f480000", x"da7c0000", x"2a230001", x"3badc9cc", x"a9b69c87", x"030a9e60", x"be0a679e", x"5fec0000", x"294b0000", x"99d20000", x"4ed00012", x"1ed34f73", x"baa708c9", x"57140bdf", x"30aebcf7"),
	(x"03790000", x"77fb0000", x"29460000", x"10e10006", x"6a84439c", x"c2d8fa98", x"0daf5183", x"58d01860", x"f7360000", x"bff50000", x"c5cf0000", x"490a0010", x"63b5daf0", x"a53f7843", x"ec7283d7", x"ea293cf7"),
	(x"a89e0000", x"e9f60000", x"86610000", x"2df90003", x"46cb5c4f", x"b62eec0d", x"b86c1668", x"648de79e", x"f40b0000", x"b7460000", x"36f50000", x"73c80017", x"329c50a0", x"ce511e5c", x"e2d74c34", x"0cf34309"),
	(x"aba30000", x"e1450000", x"755b0000", x"173b0004", x"17e2d61f", x"dd408a12", x"b6c9d98b", x"82579860", x"5cd10000", x"21f80000", x"6ae80000", x"74120015", x"4ffac523", x"d1c96ed6", x"59b1c43c", x"d674c309"),
	(x"01d70000", x"98ca0000", x"37870000", x"e52f000a", x"b67d4494", x"151528a9", x"053cff81", x"ed65f9e5", x"cdc40000", x"f5ce0000", x"ce280000", x"180c0011", x"a43a6c65", x"e048abc5", x"c7dafc8d", x"4bb8c920"),
	(x"02ea0000", x"90790000", x"c4bd0000", x"dfed000d", x"e754cec4", x"7e7b4eb6", x"0b993062", x"0bbf861b", x"651e0000", x"63700000", x"92350000", x"1fd60013", x"d95cf9e6", x"ffd0db4f", x"7cbc7485", x"913f4920"),
	(x"a90d0000", x"0e740000", x"6b9a0000", x"e2f50008", x"cb1bd117", x"0a8d5823", x"be5a7789", x"37e279e5", x"66230000", x"6bc30000", x"610f0000", x"25140014", x"887573b6", x"94bebd50", x"7219bb66", x"77e536de"),
	(x"aa300000", x"06c70000", x"98a00000", x"d837000f", x"9a325b47", x"61e33e3c", x"b0ffb86a", x"d138061b", x"cef90000", x"fd7d0000", x"3d120000", x"22ce0016", x"f513e635", x"8b26cdda", x"c97f336e", x"ad62b6de"),
	(x"926c0000", x"a3cd0000", x"8d860000", x"7cff0002", x"8144eada", x"f3593f8b", x"93c46932", x"c51c1249", x"cc570000", x"124c0000", x"23d30000", x"d700001a", x"29eae13d", x"5ceb1feb", x"c1ec9d6c", x"18d7575b"),
	(x"91510000", x"ab7e0000", x"7ebc0000", x"463d0005", x"d06d608a", x"98375994", x"9d61a6d1", x"23c66db7", x"648d0000", x"84f20000", x"7fce0000", x"d0da0018", x"548c74be", x"43736f61", x"7a8a1564", x"c250d75b"),
	(x"3ab60000", x"35730000", x"d19b0000", x"7b250000", x"fc227f59", x"ecc14f01", x"28a2e13a", x"1f9b9249", x"67b00000", x"8c410000", x"8cf40000", x"ea18001f", x"05a5feee", x"281d097e", x"742fda87", x"248aa8a5"),
	(x"398b0000", x"3dc00000", x"22a10000", x"41e70007", x"ad0bf509", x"87af291e", x"26072ed9", x"f941edb7", x"cf6a0000", x"1aff0000", x"d0e90000", x"edc2001d", x"78c36b6d", x"378579f4", x"cf49528f", x"fe0d28a5"),
	(x"93ff0000", x"444f0000", x"607d0000", x"b3f30009", x"0c946782", x"4ffa8ba5", x"95f208d3", x"96738c32", x"5e7f0000", x"cec90000", x"74290000", x"81dc0019", x"9303c22b", x"0604bce7", x"51226a3e", x"63c1228c"),
	(x"90c20000", x"4cfc0000", x"93470000", x"8931000e", x"5dbdedd2", x"2494edba", x"9b57c730", x"70a9f3cc", x"f6a50000", x"58770000", x"28340000", x"8606001b", x"ee6557a8", x"199ccc6d", x"ea44e236", x"b946a28c"),
	(x"3b250000", x"d2f10000", x"3c600000", x"b429000b", x"71f2f201", x"5062fb2f", x"2e9480db", x"4cf40c32", x"f5980000", x"50c40000", x"db0e0000", x"bcc4001c", x"bf4cddf8", x"72f2aa72", x"e4e12dd5", x"5f9cdd72"),
	(x"38180000", x"da420000", x"cf5a0000", x"8eeb000c", x"20db7851", x"3b0c9d30", x"20314f38", x"aa2e73cc", x"5d420000", x"c67a0000", x"87130000", x"bb1e001e", x"c22a487b", x"6d6adaf8", x"5f87a5dd", x"851b5d72"),
	(x"5fec0000", x"294b0000", x"99d20000", x"4ed00012", x"1ed34f73", x"baa708c9", x"57140bdf", x"30aebcf7", x"5fa80000", x"56030000", x"43ae0000", x"64f30013", x"257e86bf", x"1311944e", x"541e95bf", x"8ea4db69"),
	(x"5cd10000", x"21f80000", x"6ae80000", x"74120015", x"4ffac523", x"d1c96ed6", x"59b1c43c", x"d674c309", x"f7720000", x"c0bd0000", x"1fb30000", x"63290011", x"5818133c", x"0c89e4c4", x"ef781db7", x"54235b69"),
	(x"f7360000", x"bff50000", x"c5cf0000", x"490a0010", x"63b5daf0", x"a53f7843", x"ec7283d7", x"ea293cf7", x"f44f0000", x"c80e0000", x"ec890000", x"59eb0016", x"0931996c", x"67e782db", x"e1ddd254", x"b2f92497"),
	(x"f40b0000", x"b7460000", x"36f50000", x"73c80017", x"329c50a0", x"ce511e5c", x"e2d74c34", x"0cf34309", x"5c950000", x"5eb00000", x"b0940000", x"5e310014", x"74570cef", x"787ff251", x"5abb5a5c", x"687ea497"),
	(x"5e7f0000", x"cec90000", x"74290000", x"81dc0019", x"9303c22b", x"0604bce7", x"51226a3e", x"63c1228c", x"cd800000", x"8a860000", x"14540000", x"322f0010", x"9f97a5a9", x"49fe3742", x"c4d062ed", x"f5b2aebe"),
	(x"5d420000", x"c67a0000", x"87130000", x"bb1e001e", x"c22a487b", x"6d6adaf8", x"5f87a5dd", x"851b5d72", x"655a0000", x"1c380000", x"48490000", x"35f50012", x"e2f1302a", x"566647c8", x"7fb6eae5", x"2f352ebe"),
	(x"f6a50000", x"58770000", x"28340000", x"8606001b", x"ee6557a8", x"199ccc6d", x"ea44e236", x"b946a28c", x"66670000", x"148b0000", x"bb730000", x"0f370015", x"b3d8ba7a", x"3d0821d7", x"71132506", x"c9ef5140"),
	(x"f5980000", x"50c40000", x"db0e0000", x"bcc4001c", x"bf4cddf8", x"72f2aa72", x"e4e12dd5", x"5f9cdd72", x"cebd0000", x"82350000", x"e76e0000", x"08ed0017", x"cebe2ff9", x"2290515d", x"ca75ad0e", x"1368d140"),
	(x"cdc40000", x"f5ce0000", x"ce280000", x"180c0011", x"a43a6c65", x"e048abc5", x"c7dafc8d", x"4bb8c920", x"cc130000", x"6d040000", x"f9af0000", x"fd23001b", x"124728f1", x"f55d836c", x"c2e6030c", x"a6dd30c5"),
	(x"cef90000", x"fd7d0000", x"3d120000", x"22ce0016", x"f513e635", x"8b26cdda", x"c97f336e", x"ad62b6de", x"64c90000", x"fbba0000", x"a5b20000", x"faf90019", x"6f21bd72", x"eac5f3e6", x"79808b04", x"7c5ab0c5"),
	(x"651e0000", x"63700000", x"92350000", x"1fd60013", x"d95cf9e6", x"ffd0db4f", x"7cbc7485", x"913f4920", x"67f40000", x"f3090000", x"56880000", x"c03b001e", x"3e083722", x"81ab95f9", x"772544e7", x"9a80cf3b"),
	(x"66230000", x"6bc30000", x"610f0000", x"25140014", x"887573b6", x"94bebd50", x"7219bb66", x"77e536de", x"cf2e0000", x"65b70000", x"0a950000", x"c7e1001c", x"436ea2a1", x"9e33e573", x"cc43ccef", x"40074f3b"),
	(x"cc570000", x"124c0000", x"23d30000", x"d700001a", x"29eae13d", x"5ceb1feb", x"c1ec9d6c", x"18d7575b", x"5e3b0000", x"b1810000", x"ae550000", x"abff0018", x"a8ae0be7", x"afb22060", x"5228f45e", x"ddcb4512"),
	(x"cf6a0000", x"1aff0000", x"d0e90000", x"edc2001d", x"78c36b6d", x"378579f4", x"cf49528f", x"fe0d28a5", x"f6e10000", x"273f0000", x"f2480000", x"ac25001a", x"d5c89e64", x"b02a50ea", x"e94e7c56", x"074cc512"),
	(x"648d0000", x"84f20000", x"7fce0000", x"d0da0018", x"548c74be", x"43736f61", x"7a8a1564", x"c250d75b", x"f5dc0000", x"2f8c0000", x"01720000", x"96e7001d", x"84e11434", x"db4436f5", x"e7ebb3b5", x"e196baec"),
	(x"67b00000", x"8c410000", x"8cf40000", x"ea18001f", x"05a5feee", x"281d097e", x"742fda87", x"248aa8a5", x"5d060000", x"b9320000", x"5d6f0000", x"913d001f", x"f98781b7", x"c4dc467f", x"5c8d3bbd", x"3b113aec"),
	(x"ee930000", x"d6070000", x"92c10000", x"2b9801e0", x"9451287c", x"3b6cfb57", x"45312374", x"201f6a64", x"7b280000", x"57420000", x"a9e50000", x"634300a0", x"9edb442f", x"6d9995bb", x"27f83b03", x"c7ff60f0"),
	(x"edae0000", x"deb40000", x"61fb0000", x"115a01e7", x"c578a22c", x"50029d48", x"4b94ec97", x"c6c5159a", x"d3f20000", x"c1fc0000", x"f5f80000", x"649900a2", x"e3bdd1ac", x"7201e531", x"9c9eb30b", x"1d78e0f0"),
	(x"46490000", x"40b90000", x"cedc0000", x"2c4201e2", x"e937bdff", x"24f48bdd", x"fe57ab7c", x"fa98ea64", x"d0cf0000", x"c94f0000", x"06c20000", x"5e5b00a5", x"b2945bfc", x"196f832e", x"923b7ce8", x"fba29f0e"),
	(x"45740000", x"480a0000", x"3de60000", x"168001e5", x"b81e37af", x"4f9aedc2", x"f0f2649f", x"1c42959a", x"78150000", x"5ff10000", x"5adf0000", x"598100a7", x"cff2ce7f", x"06f7f3a4", x"295df4e0", x"21251f0e"),
	(x"ef000000", x"31850000", x"7f3a0000", x"e49401eb", x"1981a524", x"87cf4f79", x"43074295", x"7370f41f", x"e9000000", x"8bc70000", x"fe1f0000", x"359f00a3", x"24326739", x"377636b7", x"b736cc51", x"bce91527"),
	(x"ec3d0000", x"39360000", x"8c000000", x"de5601ec", x"48a82f74", x"eca12966", x"4da28d76", x"95aa8be1", x"41da0000", x"1d790000", x"a2020000", x"324500a1", x"5954f2ba", x"28ee463d", x"0c504459", x"666e9527"),
	(x"47da0000", x"a73b0000", x"23270000", x"e34e01e9", x"64e730a7", x"98573ff3", x"f861ca9d", x"a9f7741f", x"42e70000", x"15ca0000", x"51380000", x"088700a6", x"087d78ea", x"43802022", x"02f58bba", x"80b4ead9"),
	(x"44e70000", x"af880000", x"d01d0000", x"d98c01ee", x"35cebaf7", x"f33959ec", x"f6c4057e", x"4f2d0be1", x"ea3d0000", x"83740000", x"0d250000", x"0f5d00a4", x"751bed69", x"5c1850a8", x"b99303b2", x"5a336ad9"),
	(x"7cbb0000", x"0a820000", x"c53b0000", x"7d4401e3", x"2eb80b6a", x"6183585b", x"d5ffd426", x"5b091fb3", x"e8930000", x"6c450000", x"13e40000", x"fa9300a8", x"a9e2ea61", x"8bd58299", x"b100adb0", x"ef868b5c"),
	(x"7f860000", x"02310000", x"36010000", x"478601e4", x"7f91813a", x"0aed3e44", x"db5a1bc5", x"bdd3604d", x"40490000", x"fafb0000", x"4ff90000", x"fd4900aa", x"d4847fe2", x"944df213", x"0a6625b8", x"35010b5c"),
	(x"d4610000", x"9c3c0000", x"99260000", x"7a9e01e1", x"53de9ee9", x"7e1b28d1", x"6e995c2e", x"818e9fb3", x"43740000", x"f2480000", x"bcc30000", x"c78b00ad", x"85adf5b2", x"ff23940c", x"04c3ea5b", x"d3db74a2"),
	(x"d75c0000", x"948f0000", x"6a1c0000", x"405c01e6", x"02f714b9", x"15754ece", x"603c93cd", x"6754e04d", x"ebae0000", x"64f60000", x"e0de0000", x"c05100af", x"f8cb6031", x"e0bbe486", x"bfa56253", x"095cf4a2"),
	(x"7d280000", x"ed000000", x"28c00000", x"b24801e8", x"a3688632", x"dd20ec75", x"d3c9b5c7", x"086681c8", x"7abb0000", x"b0c00000", x"441e0000", x"ac4f00ab", x"130bc977", x"d13a2195", x"21ce5ae2", x"9490fe8b"),
	(x"7e150000", x"e5b30000", x"dbfa0000", x"888a01ef", x"f2410c62", x"b64e8a6a", x"dd6c7a24", x"eebcfe36", x"d2610000", x"267e0000", x"18030000", x"ab9500a9", x"6e6d5cf4", x"cea2511f", x"9aa8d2ea", x"4e177e8b"),
	(x"d5f20000", x"7bbe0000", x"74dd0000", x"b59201ea", x"de0e13b1", x"c2b89cff", x"68af3dcf", x"d2e101c8", x"d15c0000", x"2ecd0000", x"eb390000", x"915700ae", x"3f44d6a4", x"a5cc3700", x"940d1d09", x"a8cd0175"),
	(x"d6cf0000", x"730d0000", x"87e70000", x"8f5001ed", x"8f2799e1", x"a9d6fae0", x"660af22c", x"343b7e36", x"79860000", x"b8730000", x"b7240000", x"968d00ac", x"42224327", x"ba54478a", x"2f6b9501", x"724a8175"),
	(x"b13b0000", x"80040000", x"d16f0000", x"4f6b01f3", x"b12faec3", x"287d6f19", x"112fb6cb", x"aebbb10d", x"7b6c0000", x"280a0000", x"73990000", x"496000a1", x"a5768de3", x"c42f093c", x"24f2a563", x"79f5076e"),
	(x"b2060000", x"88b70000", x"22550000", x"75a901f4", x"e0062493", x"43130906", x"1f8a7928", x"4861cef3", x"d3b60000", x"beb40000", x"2f840000", x"4eba00a3", x"d8101860", x"dbb779b6", x"9f942d6b", x"a372876e"),
	(x"19e10000", x"16ba0000", x"8d720000", x"48b101f1", x"cc493b40", x"37e51f93", x"aa493ec3", x"743c310d", x"d08b0000", x"b6070000", x"dcbe0000", x"747800a4", x"89399230", x"b0d91fa9", x"9131e288", x"45a8f890"),
	(x"1adc0000", x"1e090000", x"7e480000", x"727301f6", x"9d60b110", x"5c8b798c", x"a4ecf120", x"92e64ef3", x"78510000", x"20b90000", x"80a30000", x"73a200a6", x"f45f07b3", x"af416f23", x"2a576a80", x"9f2f7890"),
	(x"b0a80000", x"67860000", x"3c940000", x"806701f8", x"3cff239b", x"94dedb37", x"1719d72a", x"fdd42f76", x"e9440000", x"f48f0000", x"24630000", x"1fbc00a2", x"1f9faef5", x"9ec0aa30", x"b43c5231", x"02e372b9"),
	(x"b3950000", x"6f350000", x"cfae0000", x"baa501ff", x"6dd6a9cb", x"ffb0bd28", x"19bc18c9", x"1b0e5088", x"419e0000", x"62310000", x"787e0000", x"186600a0", x"62f93b76", x"8158daba", x"0f5ada39", x"d864f2b9"),
	(x"18720000", x"f1380000", x"60890000", x"87bd01fa", x"4199b618", x"8b46abbd", x"ac7f5f22", x"2753af76", x"42a30000", x"6a820000", x"8b440000", x"22a400a7", x"33d0b126", x"ea36bca5", x"01ff15da", x"3ebe8d47"),
	(x"1b4f0000", x"f98b0000", x"93b30000", x"bd7f01fd", x"10b03c48", x"e028cda2", x"a2da90c1", x"c189d088", x"ea790000", x"fc3c0000", x"d7590000", x"257e00a5", x"4eb624a5", x"f5aecc2f", x"ba999dd2", x"e4390d47"),
	(x"23130000", x"5c810000", x"86950000", x"19b701f0", x"0bc68dd5", x"7292cc15", x"81e14199", x"d5adc4da", x"e8d70000", x"130d0000", x"c9980000", x"d0b000a9", x"924f23ad", x"22631e1e", x"b20a33d0", x"518cecc2"),
	(x"202e0000", x"54320000", x"75af0000", x"237501f7", x"5aef0785", x"19fcaa0a", x"8f448e7a", x"3377bb24", x"400d0000", x"85b30000", x"95850000", x"d76a00ab", x"ef29b62e", x"3dfb6e94", x"096cbbd8", x"8b0b6cc2"),
	(x"8bc90000", x"ca3f0000", x"da880000", x"1e6d01f2", x"76a01856", x"6d0abc9f", x"3a87c991", x"0f2a44da", x"43300000", x"8d000000", x"66bf0000", x"eda800ac", x"be003c7e", x"5695088b", x"07c9743b", x"6dd1133c"),
	(x"88f40000", x"c28c0000", x"29b20000", x"24af01f5", x"27899206", x"0664da80", x"34220672", x"e9f03b24", x"ebea0000", x"1bbe0000", x"3aa20000", x"ea7200ae", x"c366a9fd", x"490d7801", x"bcaffc33", x"b756933c"),
	(x"22800000", x"bb030000", x"6b6e0000", x"d6bb01fb", x"8616008d", x"ce31783b", x"87d72078", x"86c25aa1", x"7aff0000", x"cf880000", x"9e620000", x"866c00aa", x"28a600bb", x"788cbd12", x"22c4c482", x"2a9a9915"),
	(x"21bd0000", x"b3b00000", x"98540000", x"ec7901fc", x"d73f8add", x"a55f1e24", x"8972ef9b", x"6018255f", x"d2250000", x"59360000", x"c27f0000", x"81b600a8", x"55c09538", x"6714cd98", x"99a24c8a", x"f01d1915"),
	(x"8a5a0000", x"2dbd0000", x"37730000", x"d16101f9", x"fb70950e", x"d1a908b1", x"3cb1a870", x"5c45daa1", x"d1180000", x"51850000", x"31450000", x"bb7400af", x"04e91f68", x"0c7aab87", x"97078369", x"16c766eb"),
	(x"89670000", x"250e0000", x"c4490000", x"eba301fe", x"aa591f5e", x"bac76eae", x"32146793", x"ba9fa55f", x"79c20000", x"c73b0000", x"6d580000", x"bcae00ad", x"798f8aeb", x"13e2db0d", x"2c610b61", x"cc40e6eb"),
	(x"eed70000", x"a94f0000", x"48bd0000", x"01bb01e1", x"affce1b0", x"92da67d0", x"463bbd14", x"9e150dfa", x"24c40000", x"7e090000", x"30370000", x"2d9300b2", x"80080b5c", x"d73e9d72", x"70ec30dc", x"f751dc07"),
	(x"edea0000", x"a1fc0000", x"bb870000", x"3b7901e6", x"fed56be0", x"f9b401cf", x"489e72f7", x"78cf7204", x"8c1e0000", x"e8b70000", x"6c2a0000", x"2a4900b0", x"fd6e9edf", x"c8a6edf8", x"cb8ab8d4", x"2dd65c07"),
	(x"460d0000", x"3ff10000", x"14a00000", x"066101e3", x"d29a7433", x"8d42175a", x"fd5d351c", x"44928dfa", x"8f230000", x"e0040000", x"9f100000", x"108b00b7", x"ac47148f", x"a3c88be7", x"c52f7737", x"cb0c23f9"),
	(x"45300000", x"37420000", x"e79a0000", x"3ca301e4", x"83b3fe63", x"e62c7145", x"f3f8faff", x"a248f204", x"27f90000", x"76ba0000", x"c30d0000", x"175100b5", x"d121810c", x"bc50fb6d", x"7e49ff3f", x"118ba3f9"),
	(x"ef440000", x"4ecd0000", x"a5460000", x"ceb701ea", x"222c6ce8", x"2e79d3fe", x"400ddcf5", x"cd7a9381", x"b6ec0000", x"a28c0000", x"67cd0000", x"7b4f00b1", x"3ae1284a", x"8dd13e7e", x"e022c78e", x"8c47a9d0"),
	(x"ec790000", x"467e0000", x"567c0000", x"f47501ed", x"7305e6b8", x"4517b5e1", x"4ea81316", x"2ba0ec7f", x"1e360000", x"34320000", x"3bd00000", x"7c9500b3", x"4787bdc9", x"92494ef4", x"5b444f86", x"56c029d0"),
	(x"479e0000", x"d8730000", x"f95b0000", x"c96d01e8", x"5f4af96b", x"31e1a374", x"fb6b54fd", x"17fd1381", x"1d0b0000", x"3c810000", x"c8ea0000", x"465700b4", x"16ae3799", x"f92728eb", x"55e18065", x"b01a562e"),
	(x"44a30000", x"d0c00000", x"0a610000", x"f3af01ef", x"0e63733b", x"5a8fc56b", x"f5ce9b1e", x"f1276c7f", x"b5d10000", x"aa3f0000", x"94f70000", x"418d00b6", x"6bc8a21a", x"e6bf5861", x"ee87086d", x"6a9dd62e"),
	(x"7cff0000", x"75ca0000", x"1f470000", x"576701e2", x"1515c2a6", x"c835c4dc", x"d6f54a46", x"e503782d", x"b77f0000", x"450e0000", x"8a360000", x"b44300ba", x"b731a512", x"31728a50", x"e614a66f", x"df2837ab"),
	(x"7fc20000", x"7d790000", x"ec7d0000", x"6da501e5", x"443c48f6", x"a35ba2c3", x"d85085a5", x"03d907d3", x"1fa50000", x"d3b00000", x"d62b0000", x"b39900b8", x"ca573091", x"2eeafada", x"5d722e67", x"05afb7ab"),
	(x"d4250000", x"e3740000", x"435a0000", x"50bd01e0", x"68735725", x"d7adb456", x"6d93c24e", x"3f84f82d", x"1c980000", x"db030000", x"25110000", x"895b00bf", x"9b7ebac1", x"45849cc5", x"53d7e184", x"e375c855"),
	(x"d7180000", x"ebc70000", x"b0600000", x"6a7f01e7", x"395add75", x"bcc3d249", x"63360dad", x"d95e87d3", x"b4420000", x"4dbd0000", x"790c0000", x"8e8100bd", x"e6182f42", x"5a1cec4f", x"e8b1698c", x"39f24855"),
	(x"7d6c0000", x"92480000", x"f2bc0000", x"986b01e9", x"98c54ffe", x"749670f2", x"d0c32ba7", x"b66ce656", x"25570000", x"998b0000", x"ddcc0000", x"e29f00b9", x"0dd88604", x"6b9d295c", x"76da513d", x"a43e427c"),
	(x"7e510000", x"9afb0000", x"01860000", x"a2a901ee", x"c9ecc5ae", x"1ff816ed", x"de66e444", x"50b699a8", x"8d8d0000", x"0f350000", x"81d10000", x"e54500bb", x"70be1387", x"740559d6", x"cdbcd935", x"7eb9c27c"),
	(x"d5b60000", x"04f60000", x"aea10000", x"9fb101eb", x"e5a3da7d", x"6b0e0078", x"6ba5a3af", x"6ceb6656", x"8eb00000", x"07860000", x"72eb0000", x"df8700bc", x"219799d7", x"1f6b3fc9", x"c31916d6", x"9863bd82"),
	(x"d68b0000", x"0c450000", x"5d9b0000", x"a57301ec", x"b48a502d", x"00606667", x"65006c4c", x"8a3119a8", x"266a0000", x"91380000", x"2ef60000", x"d85d00be", x"5cf10c54", x"00f34f43", x"787f9ede", x"42e43d82"),
	(x"b17f0000", x"ff4c0000", x"0b130000", x"654801f2", x"8a82670f", x"81cbf39e", x"122528ab", x"10b1d693", x"24800000", x"01410000", x"ea4b0000", x"07b000b3", x"bba5c290", x"7e8801f5", x"73e6aebc", x"495bbb99"),
	(x"b2420000", x"f7ff0000", x"f8290000", x"5f8a01f5", x"dbabed5f", x"eaa59581", x"1c80e748", x"f66ba96d", x"8c5a0000", x"97ff0000", x"b6560000", x"006a00b1", x"c6c35713", x"6110717f", x"c88026b4", x"93dc3b99"),
	(x"19a50000", x"69f20000", x"570e0000", x"629201f0", x"f7e4f28c", x"9e538314", x"a943a0a3", x"ca365693", x"8f670000", x"9f4c0000", x"456c0000", x"3aa800b6", x"97eadd43", x"0a7e1760", x"c625e957", x"75064467"),
	(x"1a980000", x"61410000", x"a4340000", x"585001f7", x"a6cd78dc", x"f53de50b", x"a7e66f40", x"2cec296d", x"27bd0000", x"09f20000", x"19710000", x"3d7200b4", x"ea8c48c0", x"15e667ea", x"7d43615f", x"af81c467"),
	(x"b0ec0000", x"18ce0000", x"e6e80000", x"aa4401f9", x"0752ea57", x"3d6847b0", x"1413494a", x"43de48e8", x"b6a80000", x"ddc40000", x"bdb10000", x"516c00b0", x"014ce186", x"2467a2f9", x"e32859ee", x"324dce4e"),
	(x"b3d10000", x"107d0000", x"15d20000", x"908601fe", x"567b6007", x"560621af", x"1ab686a9", x"a5043716", x"1e720000", x"4b7a0000", x"e1ac0000", x"56b600b2", x"7c2a7405", x"3bffd273", x"584ed1e6", x"e8ca4e4e"),
	(x"18360000", x"8e700000", x"baf50000", x"ad9e01fb", x"7a347fd4", x"22f0373a", x"af75c142", x"9959c8e8", x"1d4f0000", x"43c90000", x"12960000", x"6c7400b5", x"2d03fe55", x"5091b46c", x"56eb1e05", x"0e1031b0"),
	(x"1b0b0000", x"86c30000", x"49cf0000", x"975c01fc", x"2b1df584", x"499e5125", x"a1d00ea1", x"7f83b716", x"b5950000", x"d5770000", x"4e8b0000", x"6bae00b7", x"50656bd6", x"4f09c4e6", x"ed8d960d", x"d497b1b0"),
	(x"23570000", x"23c90000", x"5ce90000", x"339401f1", x"306b4419", x"db245092", x"82ebdff9", x"6ba7a344", x"b73b0000", x"3a460000", x"504a0000", x"9e6000bb", x"8c9c6cde", x"98c416d7", x"e51e380f", x"61225035"),
	(x"206a0000", x"2b7a0000", x"afd30000", x"095601f6", x"6142ce49", x"b04a368d", x"8c4e101a", x"8d7ddcba", x"1fe10000", x"acf80000", x"0c570000", x"99ba00b9", x"f1faf95d", x"875c665d", x"5e78b007", x"bba5d035"),
	(x"8b8d0000", x"b5770000", x"00f40000", x"344e01f3", x"4d0dd19a", x"c4bc2018", x"398d57f1", x"b1202344", x"1cdc0000", x"a44b0000", x"ff6d0000", x"a37800be", x"a0d3730d", x"ec320042", x"50dd7fe4", x"5d7fafcb"),
	(x"88b00000", x"bdc40000", x"f3ce0000", x"0e8c01f4", x"1c245bca", x"afd24607", x"37289812", x"57fa5cba", x"b4060000", x"32f50000", x"a3700000", x"a4a200bc", x"ddb5e68e", x"f3aa70c8", x"ebbbf7ec", x"87f82fcb"),
	(x"22c40000", x"c44b0000", x"b1120000", x"fc9801fa", x"bdbbc941", x"6787e4bc", x"84ddbe18", x"38c83d3f", x"25130000", x"e6c30000", x"07b00000", x"c8bc00b8", x"36754fc8", x"c22bb5db", x"75d0cf5d", x"1a3425e2"),
	(x"21f90000", x"ccf80000", x"42280000", x"c65a01fd", x"ec924311", x"0ce982a3", x"8a7871fb", x"de1242c1", x"8dc90000", x"707d0000", x"5bad0000", x"cf6600ba", x"4b13da4b", x"ddb3c551", x"ceb64755", x"c0b3a5e2"),
	(x"8a1e0000", x"52f50000", x"ed0f0000", x"fb4201f8", x"c0dd5cc2", x"781f9436", x"3fbb3610", x"e24fbd3f", x"8ef40000", x"78ce0000", x"a8970000", x"f5a400bd", x"1a3a501b", x"b6dda34e", x"c01388b6", x"2669da1c"),
	(x"89230000", x"5a460000", x"1e350000", x"c18001ff", x"91f4d692", x"1371f229", x"311ef9f3", x"0495c2c1", x"262e0000", x"ee700000", x"f48a0000", x"f27e00bf", x"675cc598", x"a945d3c4", x"7b7500be", x"fcee5a1c"),
	(x"7b280000", x"57420000", x"a9e50000", x"634300a0", x"9edb442f", x"6d9995bb", x"27f83b03", x"c7ff60f0", x"95bb0000", x"81450000", x"3b240000", x"48db0140", x"0a8a6c53", x"56f56eec", x"62c91877", x"e7e00a94"),
	(x"78150000", x"5ff10000", x"5adf0000", x"598100a7", x"cff2ce7f", x"06f7f3a4", x"295df4e0", x"21251f0e", x"3d610000", x"17fb0000", x"67390000", x"4f010142", x"77ecf9d0", x"496d1e66", x"d9af907f", x"3d678a94"),
	(x"d3f20000", x"c1fc0000", x"f5f80000", x"649900a2", x"e3bdd1ac", x"7201e531", x"9c9eb30b", x"1d78e0f0", x"3e5c0000", x"1f480000", x"94030000", x"75c30145", x"26c57380", x"22037879", x"d70a5f9c", x"dbbdf56a"),
	(x"d0cf0000", x"c94f0000", x"06c20000", x"5e5b00a5", x"b2945bfc", x"196f832e", x"923b7ce8", x"fba29f0e", x"96860000", x"89f60000", x"c81e0000", x"72190147", x"5ba3e603", x"3d9b08f3", x"6c6cd794", x"013a756a"),
	(x"7abb0000", x"b0c00000", x"441e0000", x"ac4f00ab", x"130bc977", x"d13a2195", x"21ce5ae2", x"9490fe8b", x"07930000", x"5dc00000", x"6cde0000", x"1e070143", x"b0634f45", x"0c1acde0", x"f207ef25", x"9cf67f43"),
	(x"79860000", x"b8730000", x"b7240000", x"968d00ac", x"42224327", x"ba54478a", x"2f6b9501", x"724a8175", x"af490000", x"cb7e0000", x"30c30000", x"19dd0141", x"cd05dac6", x"1382bd6a", x"4961672d", x"4671ff43"),
	(x"d2610000", x"267e0000", x"18030000", x"ab9500a9", x"6e6d5cf4", x"cea2511f", x"9aa8d2ea", x"4e177e8b", x"ac740000", x"c3cd0000", x"c3f90000", x"231f0146", x"9c2c5096", x"78ecdb75", x"47c4a8ce", x"a0ab80bd"),
	(x"d15c0000", x"2ecd0000", x"eb390000", x"915700ae", x"3f44d6a4", x"a5cc3700", x"940d1d09", x"a8cd0175", x"04ae0000", x"55730000", x"9fe40000", x"24c50144", x"e14ac515", x"6774abff", x"fca220c6", x"7a2c00bd"),
	(x"e9000000", x"8bc70000", x"fe1f0000", x"359f00a3", x"24326739", x"377636b7", x"b736cc51", x"bce91527", x"06000000", x"ba420000", x"81250000", x"d10b0148", x"3db3c21d", x"b0b979ce", x"f4318ec4", x"cf99e138"),
	(x"ea3d0000", x"83740000", x"0d250000", x"0f5d00a4", x"751bed69", x"5c1850a8", x"b99303b2", x"5a336ad9", x"aeda0000", x"2cfc0000", x"dd380000", x"d6d1014a", x"40d5579e", x"af210944", x"4f5706cc", x"151e6138"),
	(x"41da0000", x"1d790000", x"a2020000", x"324500a1", x"5954f2ba", x"28ee463d", x"0c504459", x"666e9527", x"ade70000", x"244f0000", x"2e020000", x"ec13014d", x"11fcddce", x"c44f6f5b", x"41f2c92f", x"f3c41ec6"),
	(x"42e70000", x"15ca0000", x"51380000", x"088700a6", x"087d78ea", x"43802022", x"02f58bba", x"80b4ead9", x"053d0000", x"b2f10000", x"721f0000", x"ebc9014f", x"6c9a484d", x"dbd71fd1", x"fa944127", x"29439ec6"),
	(x"e8930000", x"6c450000", x"13e40000", x"fa9300a8", x"a9e2ea61", x"8bd58299", x"b100adb0", x"ef868b5c", x"94280000", x"66c70000", x"d6df0000", x"87d7014b", x"875ae10b", x"ea56dac2", x"64ff7996", x"b48f94ef"),
	(x"ebae0000", x"64f60000", x"e0de0000", x"c05100af", x"f8cb6031", x"e0bbe486", x"bfa56253", x"095cf4a2", x"3cf20000", x"f0790000", x"8ac20000", x"800d0149", x"fa3c7488", x"f5ceaa48", x"df99f19e", x"6e0814ef"),
	(x"40490000", x"fafb0000", x"4ff90000", x"fd4900aa", x"d4847fe2", x"944df213", x"0a6625b8", x"35010b5c", x"3fcf0000", x"f8ca0000", x"79f80000", x"bacf014e", x"ab15fed8", x"9ea0cc57", x"d13c3e7d", x"88d26b11"),
	(x"43740000", x"f2480000", x"bcc30000", x"c78b00ad", x"85adf5b2", x"ff23940c", x"04c3ea5b", x"d3db74a2", x"97150000", x"6e740000", x"25e50000", x"bd15014c", x"d6736b5b", x"8138bcdd", x"6a5ab675", x"5255eb11"),
	(x"24800000", x"01410000", x"ea4b0000", x"07b000b3", x"bba5c290", x"7e8801f5", x"73e6aebc", x"495bbb99", x"95ff0000", x"fe0d0000", x"e1580000", x"62f80141", x"3127a59f", x"ff43f26b", x"61c38617", x"59ea6d0a"),
	(x"27bd0000", x"09f20000", x"19710000", x"3d7200b4", x"ea8c48c0", x"15e667ea", x"7d43615f", x"af81c467", x"3d250000", x"68b30000", x"bd450000", x"65220143", x"4c41301c", x"e0db82e1", x"daa50e1f", x"836ded0a"),
	(x"8c5a0000", x"97ff0000", x"b6560000", x"006a00b1", x"c6c35713", x"6110717f", x"c88026b4", x"93dc3b99", x"3e180000", x"60000000", x"4e7f0000", x"5fe00144", x"1d68ba4c", x"8bb5e4fe", x"d400c1fc", x"65b792f4"),
	(x"8f670000", x"9f4c0000", x"456c0000", x"3aa800b6", x"97eadd43", x"0a7e1760", x"c625e957", x"75064467", x"96c20000", x"f6be0000", x"12620000", x"583a0146", x"600e2fcf", x"942d9474", x"6f6649f4", x"bf3012f4"),
	(x"25130000", x"e6c30000", x"07b00000", x"c8bc00b8", x"36754fc8", x"c22bb5db", x"75d0cf5d", x"1a3425e2", x"07d70000", x"22880000", x"b6a20000", x"34240142", x"8bce8689", x"a5ac5167", x"f10d7145", x"22fc18dd"),
	(x"262e0000", x"ee700000", x"f48a0000", x"f27e00bf", x"675cc598", x"a945d3c4", x"7b7500be", x"fcee5a1c", x"af0d0000", x"b4360000", x"eabf0000", x"33fe0140", x"f6a8130a", x"ba3421ed", x"4a6bf94d", x"f87b98dd"),
	(x"8dc90000", x"707d0000", x"5bad0000", x"cf6600ba", x"4b13da4b", x"ddb3c551", x"ceb64755", x"c0b3a5e2", x"ac300000", x"bc850000", x"19850000", x"093c0147", x"a781995a", x"d15a47f2", x"44ce36ae", x"1ea1e723"),
	(x"8ef40000", x"78ce0000", x"a8970000", x"f5a400bd", x"1a3a501b", x"b6dda34e", x"c01388b6", x"2669da1c", x"04ea0000", x"2a3b0000", x"45980000", x"0ee60145", x"dae70cd9", x"cec23778", x"ffa8bea6", x"c4266723"),
	(x"b6a80000", x"ddc40000", x"bdb10000", x"516c00b0", x"014ce186", x"2467a2f9", x"e32859ee", x"324dce4e", x"06440000", x"c50a0000", x"5b590000", x"fb280149", x"061e0bd1", x"190fe549", x"f73b10a4", x"719386a6"),
	(x"b5950000", x"d5770000", x"4e8b0000", x"6bae00b7", x"50656bd6", x"4f09c4e6", x"ed8d960d", x"d497b1b0", x"ae9e0000", x"53b40000", x"07440000", x"fcf2014b", x"7b789e52", x"069795c3", x"4c5d98ac", x"ab1406a6"),
	(x"1e720000", x"4b7a0000", x"e1ac0000", x"56b600b2", x"7c2a7405", x"3bffd273", x"584ed1e6", x"e8ca4e4e", x"ada30000", x"5b070000", x"f47e0000", x"c630014c", x"2a511402", x"6df9f3dc", x"42f8574f", x"4dce7958"),
	(x"1d4f0000", x"43c90000", x"12960000", x"6c7400b5", x"2d03fe55", x"5091b46c", x"56eb1e05", x"0e1031b0", x"05790000", x"cdb90000", x"a8630000", x"c1ea014e", x"57378181", x"72618356", x"f99edf47", x"9749f958"),
	(x"b73b0000", x"3a460000", x"504a0000", x"9e6000bb", x"8c9c6cde", x"98c416d7", x"e51e380f", x"61225035", x"946c0000", x"198f0000", x"0ca30000", x"adf4014a", x"bcf728c7", x"43e04645", x"67f5e7f6", x"0a85f371"),
	(x"b4060000", x"32f50000", x"a3700000", x"a4a200bc", x"ddb5e68e", x"f3aa70c8", x"ebbbf7ec", x"87f82fcb", x"3cb60000", x"8f310000", x"50be0000", x"aa2e0148", x"c191bd44", x"5c7836cf", x"dc936ffe", x"d0027371"),
	(x"1fe10000", x"acf80000", x"0c570000", x"99ba00b9", x"f1faf95d", x"875c665d", x"5e78b007", x"bba5d035", x"3f8b0000", x"87820000", x"a3840000", x"90ec014f", x"90b83714", x"371650d0", x"d236a01d", x"36d80c8f"),
	(x"1cdc0000", x"a44b0000", x"ff6d0000", x"a37800be", x"a0d3730d", x"ec320042", x"50dd7fe4", x"5d7fafcb", x"97510000", x"113c0000", x"ff990000", x"9736014d", x"eddea297", x"288e205a", x"69502815", x"ec5f8c8f"),
	(x"7b6c0000", x"280a0000", x"73990000", x"496000a1", x"a5768de3", x"c42f093c", x"24f2a563", x"79f5076e", x"ca570000", x"a80e0000", x"a2f60000", x"060b0152", x"14592320", x"ec526625", x"35dd13a8", x"d74eb663"),
	(x"78510000", x"20b90000", x"80a30000", x"73a200a6", x"f45f07b3", x"af416f23", x"2a576a80", x"9f2f7890", x"628d0000", x"3eb00000", x"feeb0000", x"01d10150", x"693fb6a3", x"f3ca16af", x"8ebb9ba0", x"0dc93663"),
	(x"d3b60000", x"beb40000", x"2f840000", x"4eba00a3", x"d8101860", x"dbb779b6", x"9f942d6b", x"a372876e", x"61b00000", x"36030000", x"0dd10000", x"3b130157", x"38163cf3", x"98a470b0", x"801e5443", x"eb13499d"),
	(x"d08b0000", x"b6070000", x"dcbe0000", x"747800a4", x"89399230", x"b0d91fa9", x"9131e288", x"45a8f890", x"c96a0000", x"a0bd0000", x"51cc0000", x"3cc90155", x"4570a970", x"873c003a", x"3b78dc4b", x"3194c99d"),
	(x"7aff0000", x"cf880000", x"9e620000", x"866c00aa", x"28a600bb", x"788cbd12", x"22c4c482", x"2a9a9915", x"587f0000", x"748b0000", x"f50c0000", x"50d70151", x"aeb00036", x"b6bdc529", x"a513e4fa", x"ac58c3b4"),
	(x"79c20000", x"c73b0000", x"6d580000", x"bcae00ad", x"798f8aeb", x"13e2db0d", x"2c610b61", x"cc40e6eb", x"f0a50000", x"e2350000", x"a9110000", x"570d0153", x"d3d695b5", x"a925b5a3", x"1e756cf2", x"76df43b4"),
	(x"d2250000", x"59360000", x"c27f0000", x"81b600a8", x"55c09538", x"6714cd98", x"99a24c8a", x"f01d1915", x"f3980000", x"ea860000", x"5a2b0000", x"6dcf0154", x"82ff1fe5", x"c24bd3bc", x"10d0a311", x"90053c4a"),
	(x"d1180000", x"51850000", x"31450000", x"bb7400af", x"04e91f68", x"0c7aab87", x"97078369", x"16c766eb", x"5b420000", x"7c380000", x"06360000", x"6a150156", x"ff998a66", x"ddd3a336", x"abb62b19", x"4a82bc4a"),
	(x"e9440000", x"f48f0000", x"24630000", x"1fbc00a2", x"1f9faef5", x"9ec0aa30", x"b43c5231", x"02e372b9", x"59ec0000", x"93090000", x"18f70000", x"9fdb015a", x"23608d6e", x"0a1e7107", x"a325851b", x"ff375dcf"),
	(x"ea790000", x"fc3c0000", x"d7590000", x"257e00a5", x"4eb624a5", x"f5aecc2f", x"ba999dd2", x"e4390d47", x"f1360000", x"05b70000", x"44ea0000", x"98010158", x"5e0618ed", x"1586018d", x"18430d13", x"25b0ddcf"),
	(x"419e0000", x"62310000", x"787e0000", x"186600a0", x"62f93b76", x"8158daba", x"0f5ada39", x"d864f2b9", x"f20b0000", x"0d040000", x"b7d00000", x"a2c3015f", x"0f2f92bd", x"7ee86792", x"16e6c2f0", x"c36aa231"),
	(x"42a30000", x"6a820000", x"8b440000", x"22a400a7", x"33d0b126", x"ea36bca5", x"01ff15da", x"3ebe8d47", x"5ad10000", x"9bba0000", x"ebcd0000", x"a519015d", x"7249073e", x"61701718", x"ad804af8", x"19ed2231"),
	(x"e8d70000", x"130d0000", x"c9980000", x"d0b000a9", x"924f23ad", x"22631e1e", x"b20a33d0", x"518cecc2", x"cbc40000", x"4f8c0000", x"4f0d0000", x"c9070159", x"9989ae78", x"50f1d20b", x"33eb7249", x"84212818"),
	(x"ebea0000", x"1bbe0000", x"3aa20000", x"ea7200ae", x"c366a9fd", x"490d7801", x"bcaffc33", x"b756933c", x"631e0000", x"d9320000", x"13100000", x"cedd015b", x"e4ef3bfb", x"4f69a281", x"888dfa41", x"5ea6a818"),
	(x"400d0000", x"85b30000", x"95850000", x"d76a00ab", x"ef29b62e", x"3dfb6e94", x"096cbbd8", x"8b0b6cc2", x"60230000", x"d1810000", x"e02a0000", x"f41f015c", x"b5c6b1ab", x"2407c49e", x"862835a2", x"b87cd7e6"),
	(x"43300000", x"8d000000", x"66bf0000", x"eda800ac", x"be003c7e", x"5695088b", x"07c9743b", x"6dd1133c", x"c8f90000", x"473f0000", x"bc370000", x"f3c5015e", x"c8a02428", x"3b9fb414", x"3d4ebdaa", x"62fb57e6"),
	(x"24c40000", x"7e090000", x"30370000", x"2d9300b2", x"80080b5c", x"d73e9d72", x"70ec30dc", x"f751dc07", x"ca130000", x"d7460000", x"788a0000", x"2c280153", x"2ff4eaec", x"45e4faa2", x"36d78dc8", x"6944d1fd"),
	(x"27f90000", x"76ba0000", x"c30d0000", x"175100b5", x"d121810c", x"bc50fb6d", x"7e49ff3f", x"118ba3f9", x"62c90000", x"41f80000", x"24970000", x"2bf20151", x"52927f6f", x"5a7c8a28", x"8db105c0", x"b3c351fd"),
	(x"8c1e0000", x"e8b70000", x"6c2a0000", x"2a4900b0", x"fd6e9edf", x"c8a6edf8", x"cb8ab8d4", x"2dd65c07", x"61f40000", x"494b0000", x"d7ad0000", x"11300156", x"03bbf53f", x"3112ec37", x"8314ca23", x"55192e03"),
	(x"8f230000", x"e0040000", x"9f100000", x"108b00b7", x"ac47148f", x"a3c88be7", x"c52f7737", x"cb0c23f9", x"c92e0000", x"dff50000", x"8bb00000", x"16ea0154", x"7edd60bc", x"2e8a9cbd", x"3872422b", x"8f9eae03"),
	(x"25570000", x"998b0000", x"ddcc0000", x"e29f00b9", x"0dd88604", x"6b9d295c", x"76da513d", x"a43e427c", x"583b0000", x"0bc30000", x"2f700000", x"7af40150", x"951dc9fa", x"1f0b59ae", x"a6197a9a", x"1252a42a"),
	(x"266a0000", x"91380000", x"2ef60000", x"d85d00be", x"5cf10c54", x"00f34f43", x"787f9ede", x"42e43d82", x"f0e10000", x"9d7d0000", x"736d0000", x"7d2e0152", x"e87b5c79", x"00932924", x"1d7ff292", x"c8d5242a"),
	(x"8d8d0000", x"0f350000", x"81d10000", x"e54500bb", x"70be1387", x"740559d6", x"cdbcd935", x"7eb9c27c", x"f3dc0000", x"95ce0000", x"80570000", x"47ec0155", x"b952d629", x"6bfd4f3b", x"13da3d71", x"2e0f5bd4"),
	(x"8eb00000", x"07860000", x"72eb0000", x"df8700bc", x"219799d7", x"1f6b3fc9", x"c31916d6", x"9863bd82", x"5b060000", x"03700000", x"dc4a0000", x"40360157", x"c43443aa", x"74653fb1", x"a8bcb579", x"f488dbd4"),
	(x"b6ec0000", x"a28c0000", x"67cd0000", x"7b4f00b1", x"3ae1284a", x"8dd13e7e", x"e022c78e", x"8c47a9d0", x"59a80000", x"ec410000", x"c28b0000", x"b5f8015b", x"18cd44a2", x"a3a8ed80", x"a02f1b7b", x"413d3a51"),
	(x"b5d10000", x"aa3f0000", x"94f70000", x"418d00b6", x"6bc8a21a", x"e6bf5861", x"ee87086d", x"6a9dd62e", x"f1720000", x"7aff0000", x"9e960000", x"b2220159", x"65abd121", x"bc309d0a", x"1b499373", x"9bbaba51"),
	(x"1e360000", x"34320000", x"3bd00000", x"7c9500b3", x"4787bdc9", x"92494ef4", x"5b444f86", x"56c029d0", x"f24f0000", x"724c0000", x"6dac0000", x"88e0015e", x"34825b71", x"d75efb15", x"15ec5c90", x"7d60c5af"),
	(x"1d0b0000", x"3c810000", x"c8ea0000", x"465700b4", x"16ae3799", x"f92728eb", x"55e18065", x"b01a562e", x"5a950000", x"e4f20000", x"31b10000", x"8f3a015c", x"49e4cef2", x"c8c68b9f", x"ae8ad498", x"a7e745af"),
	(x"b77f0000", x"450e0000", x"8a360000", x"b44300ba", x"b731a512", x"31728a50", x"e614a66f", x"df2837ab", x"cb800000", x"30c40000", x"95710000", x"e3240158", x"a22467b4", x"f9474e8c", x"30e1ec29", x"3a2b4f86"),
	(x"b4420000", x"4dbd0000", x"790c0000", x"8e8100bd", x"e6182f42", x"5a1cec4f", x"e8b1698c", x"39f24855", x"635a0000", x"a67a0000", x"c96c0000", x"e4fe015a", x"df42f237", x"e6df3e06", x"8b876421", x"e0accf86"),
	(x"1fa50000", x"d3b00000", x"d62b0000", x"b39900b8", x"ca573091", x"2eeafada", x"5d722e67", x"05afb7ab", x"60670000", x"aec90000", x"3a560000", x"de3c015d", x"8e6b7867", x"8db15819", x"8522abc2", x"0676b078"),
	(x"1c980000", x"db030000", x"25110000", x"895b00bf", x"9b7ebac1", x"45849cc5", x"53d7e184", x"e375c855", x"c8bd0000", x"38770000", x"664b0000", x"d9e6015f", x"f30dede4", x"92292893", x"3e4423ca", x"dcf13078"),
	(x"95bb0000", x"81450000", x"3b240000", x"48db0140", x"0a8a6c53", x"56f56eec", x"62c91877", x"e7e00a94", x"ee930000", x"d6070000", x"92c10000", x"2b9801e0", x"9451287c", x"3b6cfb57", x"45312374", x"201f6a64"),
	(x"96860000", x"89f60000", x"c81e0000", x"72190147", x"5ba3e603", x"3d9b08f3", x"6c6cd794", x"013a756a", x"46490000", x"40b90000", x"cedc0000", x"2c4201e2", x"e937bdff", x"24f48bdd", x"fe57ab7c", x"fa98ea64"),
	(x"3d610000", x"17fb0000", x"67390000", x"4f010142", x"77ecf9d0", x"496d1e66", x"d9af907f", x"3d678a94", x"45740000", x"480a0000", x"3de60000", x"168001e5", x"b81e37af", x"4f9aedc2", x"f0f2649f", x"1c42959a"),
	(x"3e5c0000", x"1f480000", x"94030000", x"75c30145", x"26c57380", x"22037879", x"d70a5f9c", x"dbbdf56a", x"edae0000", x"deb40000", x"61fb0000", x"115a01e7", x"c578a22c", x"50029d48", x"4b94ec97", x"c6c5159a"),
	(x"94280000", x"66c70000", x"d6df0000", x"87d7014b", x"875ae10b", x"ea56dac2", x"64ff7996", x"b48f94ef", x"7cbb0000", x"0a820000", x"c53b0000", x"7d4401e3", x"2eb80b6a", x"6183585b", x"d5ffd426", x"5b091fb3"),
	(x"97150000", x"6e740000", x"25e50000", x"bd15014c", x"d6736b5b", x"8138bcdd", x"6a5ab675", x"5255eb11", x"d4610000", x"9c3c0000", x"99260000", x"7a9e01e1", x"53de9ee9", x"7e1b28d1", x"6e995c2e", x"818e9fb3"),
	(x"3cf20000", x"f0790000", x"8ac20000", x"800d0149", x"fa3c7488", x"f5ceaa48", x"df99f19e", x"6e0814ef", x"d75c0000", x"948f0000", x"6a1c0000", x"405c01e6", x"02f714b9", x"15754ece", x"603c93cd", x"6754e04d"),
	(x"3fcf0000", x"f8ca0000", x"79f80000", x"bacf014e", x"ab15fed8", x"9ea0cc57", x"d13c3e7d", x"88d26b11", x"7f860000", x"02310000", x"36010000", x"478601e4", x"7f91813a", x"0aed3e44", x"db5a1bc5", x"bdd3604d"),
	(x"07930000", x"5dc00000", x"6cde0000", x"1e070143", x"b0634f45", x"0c1acde0", x"f207ef25", x"9cf67f43", x"7d280000", x"ed000000", x"28c00000", x"b24801e8", x"a3688632", x"dd20ec75", x"d3c9b5c7", x"086681c8"),
	(x"04ae0000", x"55730000", x"9fe40000", x"24c50144", x"e14ac515", x"6774abff", x"fca220c6", x"7a2c00bd", x"d5f20000", x"7bbe0000", x"74dd0000", x"b59201ea", x"de0e13b1", x"c2b89cff", x"68af3dcf", x"d2e101c8"),
	(x"af490000", x"cb7e0000", x"30c30000", x"19dd0141", x"cd05dac6", x"1382bd6a", x"4961672d", x"4671ff43", x"d6cf0000", x"730d0000", x"87e70000", x"8f5001ed", x"8f2799e1", x"a9d6fae0", x"660af22c", x"343b7e36"),
	(x"ac740000", x"c3cd0000", x"c3f90000", x"231f0146", x"9c2c5096", x"78ecdb75", x"47c4a8ce", x"a0ab80bd", x"7e150000", x"e5b30000", x"dbfa0000", x"888a01ef", x"f2410c62", x"b64e8a6a", x"dd6c7a24", x"eebcfe36"),
	(x"06000000", x"ba420000", x"81250000", x"d10b0148", x"3db3c21d", x"b0b979ce", x"f4318ec4", x"cf99e138", x"ef000000", x"31850000", x"7f3a0000", x"e49401eb", x"1981a524", x"87cf4f79", x"43074295", x"7370f41f"),
	(x"053d0000", x"b2f10000", x"721f0000", x"ebc9014f", x"6c9a484d", x"dbd71fd1", x"fa944127", x"29439ec6", x"47da0000", x"a73b0000", x"23270000", x"e34e01e9", x"64e730a7", x"98573ff3", x"f861ca9d", x"a9f7741f"),
	(x"aeda0000", x"2cfc0000", x"dd380000", x"d6d1014a", x"40d5579e", x"af210944", x"4f5706cc", x"151e6138", x"44e70000", x"af880000", x"d01d0000", x"d98c01ee", x"35cebaf7", x"f33959ec", x"f6c4057e", x"4f2d0be1"),
	(x"ade70000", x"244f0000", x"2e020000", x"ec13014d", x"11fcddce", x"c44f6f5b", x"41f2c92f", x"f3c41ec6", x"ec3d0000", x"39360000", x"8c000000", x"de5601ec", x"48a82f74", x"eca12966", x"4da28d76", x"95aa8be1"),
	(x"ca130000", x"d7460000", x"788a0000", x"2c280153", x"2ff4eaec", x"45e4faa2", x"36d78dc8", x"6944d1fd", x"eed70000", x"a94f0000", x"48bd0000", x"01bb01e1", x"affce1b0", x"92da67d0", x"463bbd14", x"9e150dfa"),
	(x"c92e0000", x"dff50000", x"8bb00000", x"16ea0154", x"7edd60bc", x"2e8a9cbd", x"3872422b", x"8f9eae03", x"460d0000", x"3ff10000", x"14a00000", x"066101e3", x"d29a7433", x"8d42175a", x"fd5d351c", x"44928dfa"),
	(x"62c90000", x"41f80000", x"24970000", x"2bf20151", x"52927f6f", x"5a7c8a28", x"8db105c0", x"b3c351fd", x"45300000", x"37420000", x"e79a0000", x"3ca301e4", x"83b3fe63", x"e62c7145", x"f3f8faff", x"a248f204"),
	(x"61f40000", x"494b0000", x"d7ad0000", x"11300156", x"03bbf53f", x"3112ec37", x"8314ca23", x"55192e03", x"edea0000", x"a1fc0000", x"bb870000", x"3b7901e6", x"fed56be0", x"f9b401cf", x"489e72f7", x"78cf7204"),
	(x"cb800000", x"30c40000", x"95710000", x"e3240158", x"a22467b4", x"f9474e8c", x"30e1ec29", x"3a2b4f86", x"7cff0000", x"75ca0000", x"1f470000", x"576701e2", x"1515c2a6", x"c835c4dc", x"d6f54a46", x"e503782d"),
	(x"c8bd0000", x"38770000", x"664b0000", x"d9e6015f", x"f30dede4", x"92292893", x"3e4423ca", x"dcf13078", x"d4250000", x"e3740000", x"435a0000", x"50bd01e0", x"68735725", x"d7adb456", x"6d93c24e", x"3f84f82d"),
	(x"635a0000", x"a67a0000", x"c96c0000", x"e4fe015a", x"df42f237", x"e6df3e06", x"8b876421", x"e0accf86", x"d7180000", x"ebc70000", x"b0600000", x"6a7f01e7", x"395add75", x"bcc3d249", x"63360dad", x"d95e87d3"),
	(x"60670000", x"aec90000", x"3a560000", x"de3c015d", x"8e6b7867", x"8db15819", x"8522abc2", x"0676b078", x"7fc20000", x"7d790000", x"ec7d0000", x"6da501e5", x"443c48f6", x"a35ba2c3", x"d85085a5", x"03d907d3"),
	(x"583b0000", x"0bc30000", x"2f700000", x"7af40150", x"951dc9fa", x"1f0b59ae", x"a6197a9a", x"1252a42a", x"7d6c0000", x"92480000", x"f2bc0000", x"986b01e9", x"98c54ffe", x"749670f2", x"d0c32ba7", x"b66ce656"),
	(x"5b060000", x"03700000", x"dc4a0000", x"40360157", x"c43443aa", x"74653fb1", x"a8bcb579", x"f488dbd4", x"d5b60000", x"04f60000", x"aea10000", x"9fb101eb", x"e5a3da7d", x"6b0e0078", x"6ba5a3af", x"6ceb6656"),
	(x"f0e10000", x"9d7d0000", x"736d0000", x"7d2e0152", x"e87b5c79", x"00932924", x"1d7ff292", x"c8d5242a", x"d68b0000", x"0c450000", x"5d9b0000", x"a57301ec", x"b48a502d", x"00606667", x"65006c4c", x"8a3119a8"),
	(x"f3dc0000", x"95ce0000", x"80570000", x"47ec0155", x"b952d629", x"6bfd4f3b", x"13da3d71", x"2e0f5bd4", x"7e510000", x"9afb0000", x"01860000", x"a2a901ee", x"c9ecc5ae", x"1ff816ed", x"de66e444", x"50b699a8"),
	(x"59a80000", x"ec410000", x"c28b0000", x"b5f8015b", x"18cd44a2", x"a3a8ed80", x"a02f1b7b", x"413d3a51", x"ef440000", x"4ecd0000", x"a5460000", x"ceb701ea", x"222c6ce8", x"2e79d3fe", x"400ddcf5", x"cd7a9381"),
	(x"5a950000", x"e4f20000", x"31b10000", x"8f3a015c", x"49e4cef2", x"c8c68b9f", x"ae8ad498", x"a7e745af", x"479e0000", x"d8730000", x"f95b0000", x"c96d01e8", x"5f4af96b", x"31e1a374", x"fb6b54fd", x"17fd1381"),
	(x"f1720000", x"7aff0000", x"9e960000", x"b2220159", x"65abd121", x"bc309d0a", x"1b499373", x"9bbaba51", x"44a30000", x"d0c00000", x"0a610000", x"f3af01ef", x"0e63733b", x"5a8fc56b", x"f5ce9b1e", x"f1276c7f"),
	(x"f24f0000", x"724c0000", x"6dac0000", x"88e0015e", x"34825b71", x"d75efb15", x"15ec5c90", x"7d60c5af", x"ec790000", x"467e0000", x"567c0000", x"f47501ed", x"7305e6b8", x"4517b5e1", x"4ea81316", x"2ba0ec7f"),
	(x"95ff0000", x"fe0d0000", x"e1580000", x"62f80141", x"3127a59f", x"ff43f26b", x"61c38617", x"59ea6d0a", x"b17f0000", x"ff4c0000", x"0b130000", x"654801f2", x"8a82670f", x"81cbf39e", x"122528ab", x"10b1d693"),
	(x"96c20000", x"f6be0000", x"12620000", x"583a0146", x"600e2fcf", x"942d9474", x"6f6649f4", x"bf3012f4", x"19a50000", x"69f20000", x"570e0000", x"629201f0", x"f7e4f28c", x"9e538314", x"a943a0a3", x"ca365693"),
	(x"3d250000", x"68b30000", x"bd450000", x"65220143", x"4c41301c", x"e0db82e1", x"daa50e1f", x"836ded0a", x"1a980000", x"61410000", x"a4340000", x"585001f7", x"a6cd78dc", x"f53de50b", x"a7e66f40", x"2cec296d"),
	(x"3e180000", x"60000000", x"4e7f0000", x"5fe00144", x"1d68ba4c", x"8bb5e4fe", x"d400c1fc", x"65b792f4", x"b2420000", x"f7ff0000", x"f8290000", x"5f8a01f5", x"dbabed5f", x"eaa59581", x"1c80e748", x"f66ba96d"),
	(x"946c0000", x"198f0000", x"0ca30000", x"adf4014a", x"bcf728c7", x"43e04645", x"67f5e7f6", x"0a85f371", x"23570000", x"23c90000", x"5ce90000", x"339401f1", x"306b4419", x"db245092", x"82ebdff9", x"6ba7a344"),
	(x"97510000", x"113c0000", x"ff990000", x"9736014d", x"eddea297", x"288e205a", x"69502815", x"ec5f8c8f", x"8b8d0000", x"b5770000", x"00f40000", x"344e01f3", x"4d0dd19a", x"c4bc2018", x"398d57f1", x"b1202344"),
	(x"3cb60000", x"8f310000", x"50be0000", x"aa2e0148", x"c191bd44", x"5c7836cf", x"dc936ffe", x"d0027371", x"88b00000", x"bdc40000", x"f3ce0000", x"0e8c01f4", x"1c245bca", x"afd24607", x"37289812", x"57fa5cba"),
	(x"3f8b0000", x"87820000", x"a3840000", x"90ec014f", x"90b83714", x"371650d0", x"d236a01d", x"36d80c8f", x"206a0000", x"2b7a0000", x"afd30000", x"095601f6", x"6142ce49", x"b04a368d", x"8c4e101a", x"8d7ddcba"),
	(x"07d70000", x"22880000", x"b6a20000", x"34240142", x"8bce8689", x"a5ac5167", x"f10d7145", x"22fc18dd", x"22c40000", x"c44b0000", x"b1120000", x"fc9801fa", x"bdbbc941", x"6787e4bc", x"84ddbe18", x"38c83d3f"),
	(x"04ea0000", x"2a3b0000", x"45980000", x"0ee60145", x"dae70cd9", x"cec23778", x"ffa8bea6", x"c4266723", x"8a1e0000", x"52f50000", x"ed0f0000", x"fb4201f8", x"c0dd5cc2", x"781f9436", x"3fbb3610", x"e24fbd3f"),
	(x"af0d0000", x"b4360000", x"eabf0000", x"33fe0140", x"f6a8130a", x"ba3421ed", x"4a6bf94d", x"f87b98dd", x"89230000", x"5a460000", x"1e350000", x"c18001ff", x"91f4d692", x"1371f229", x"311ef9f3", x"0495c2c1"),
	(x"ac300000", x"bc850000", x"19850000", x"093c0147", x"a781995a", x"d15a47f2", x"44ce36ae", x"1ea1e723", x"21f90000", x"ccf80000", x"42280000", x"c65a01fd", x"ec924311", x"0ce982a3", x"8a7871fb", x"de1242c1"),
	(x"06440000", x"c50a0000", x"5b590000", x"fb280149", x"061e0bd1", x"190fe549", x"f73b10a4", x"719386a6", x"b0ec0000", x"18ce0000", x"e6e80000", x"aa4401f9", x"0752ea57", x"3d6847b0", x"1413494a", x"43de48e8"),
	(x"05790000", x"cdb90000", x"a8630000", x"c1ea014e", x"57378181", x"72618356", x"f99edf47", x"9749f958", x"18360000", x"8e700000", x"baf50000", x"ad9e01fb", x"7a347fd4", x"22f0373a", x"af75c142", x"9959c8e8"),
	(x"ae9e0000", x"53b40000", x"07440000", x"fcf2014b", x"7b789e52", x"069795c3", x"4c5d98ac", x"ab1406a6", x"1b0b0000", x"86c30000", x"49cf0000", x"975c01fc", x"2b1df584", x"499e5125", x"a1d00ea1", x"7f83b716"),
	(x"ada30000", x"5b070000", x"f47e0000", x"c630014c", x"2a511402", x"6df9f3dc", x"42f8574f", x"4dce7958", x"b3d10000", x"107d0000", x"15d20000", x"908601fe", x"567b6007", x"560621af", x"1ab686a9", x"a5043716"),
	(x"ca570000", x"a80e0000", x"a2f60000", x"060b0152", x"14592320", x"ec526625", x"35dd13a8", x"d74eb663", x"b13b0000", x"80040000", x"d16f0000", x"4f6b01f3", x"b12faec3", x"287d6f19", x"112fb6cb", x"aebbb10d"),
	(x"c96a0000", x"a0bd0000", x"51cc0000", x"3cc90155", x"4570a970", x"873c003a", x"3b78dc4b", x"3194c99d", x"19e10000", x"16ba0000", x"8d720000", x"48b101f1", x"cc493b40", x"37e51f93", x"aa493ec3", x"743c310d"),
	(x"628d0000", x"3eb00000", x"feeb0000", x"01d10150", x"693fb6a3", x"f3ca16af", x"8ebb9ba0", x"0dc93663", x"1adc0000", x"1e090000", x"7e480000", x"727301f6", x"9d60b110", x"5c8b798c", x"a4ecf120", x"92e64ef3"),
	(x"61b00000", x"36030000", x"0dd10000", x"3b130157", x"38163cf3", x"98a470b0", x"801e5443", x"eb13499d", x"b2060000", x"88b70000", x"22550000", x"75a901f4", x"e0062493", x"43130906", x"1f8a7928", x"4861cef3"),
	(x"cbc40000", x"4f8c0000", x"4f0d0000", x"c9070159", x"9989ae78", x"50f1d20b", x"33eb7249", x"84212818", x"23130000", x"5c810000", x"86950000", x"19b701f0", x"0bc68dd5", x"7292cc15", x"81e14199", x"d5adc4da"),
	(x"c8f90000", x"473f0000", x"bc370000", x"f3c5015e", x"c8a02428", x"3b9fb414", x"3d4ebdaa", x"62fb57e6", x"8bc90000", x"ca3f0000", x"da880000", x"1e6d01f2", x"76a01856", x"6d0abc9f", x"3a87c991", x"0f2a44da"),
	(x"631e0000", x"d9320000", x"13100000", x"cedd015b", x"e4ef3bfb", x"4f69a281", x"888dfa41", x"5ea6a818", x"88f40000", x"c28c0000", x"29b20000", x"24af01f5", x"27899206", x"0664da80", x"34220672", x"e9f03b24"),
	(x"60230000", x"d1810000", x"e02a0000", x"f41f015c", x"b5c6b1ab", x"2407c49e", x"862835a2", x"b87cd7e6", x"202e0000", x"54320000", x"75af0000", x"237501f7", x"5aef0785", x"19fcaa0a", x"8f448e7a", x"3377bb24"),
	(x"587f0000", x"748b0000", x"f50c0000", x"50d70151", x"aeb00036", x"b6bdc529", x"a513e4fa", x"ac58c3b4", x"22800000", x"bb030000", x"6b6e0000", x"d6bb01fb", x"8616008d", x"ce31783b", x"87d72078", x"86c25aa1"),
	(x"5b420000", x"7c380000", x"06360000", x"6a150156", x"ff998a66", x"ddd3a336", x"abb62b19", x"4a82bc4a", x"8a5a0000", x"2dbd0000", x"37730000", x"d16101f9", x"fb70950e", x"d1a908b1", x"3cb1a870", x"5c45daa1"),
	(x"f0a50000", x"e2350000", x"a9110000", x"570d0153", x"d3d695b5", x"a925b5a3", x"1e756cf2", x"76df43b4", x"89670000", x"250e0000", x"c4490000", x"eba301fe", x"aa591f5e", x"bac76eae", x"32146793", x"ba9fa55f"),
	(x"f3980000", x"ea860000", x"5a2b0000", x"6dcf0154", x"82ff1fe5", x"c24bd3bc", x"10d0a311", x"90053c4a", x"21bd0000", x"b3b00000", x"98540000", x"ec7901fc", x"d73f8add", x"a55f1e24", x"8972ef9b", x"6018255f"),
	(x"59ec0000", x"93090000", x"18f70000", x"9fdb015a", x"23608d6e", x"0a1e7107", x"a325851b", x"ff375dcf", x"b0a80000", x"67860000", x"3c940000", x"806701f8", x"3cff239b", x"94dedb37", x"1719d72a", x"fdd42f76"),
	(x"5ad10000", x"9bba0000", x"ebcd0000", x"a519015d", x"7249073e", x"61701718", x"ad804af8", x"19ed2231", x"18720000", x"f1380000", x"60890000", x"87bd01fa", x"4199b618", x"8b46abbd", x"ac7f5f22", x"2753af76"),
	(x"f1360000", x"05b70000", x"44ea0000", x"98010158", x"5e0618ed", x"1586018d", x"18430d13", x"25b0ddcf", x"1b4f0000", x"f98b0000", x"93b30000", x"bd7f01fd", x"10b03c48", x"e028cda2", x"a2da90c1", x"c189d088"),
	(x"f20b0000", x"0d040000", x"b7d00000", x"a2c3015f", x"0f2f92bd", x"7ee86792", x"16e6c2f0", x"c36aa231", x"b3950000", x"6f350000", x"cfae0000", x"baa501ff", x"6dd6a9cb", x"ffb0bd28", x"19bc18c9", x"1b0e5088")
    ));

	
end package;