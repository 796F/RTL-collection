-- =====================================================================
-- Copyright � 2010 by Cryptographic Engineering Research Group (CERG),
-- ECE Department, George Mason University
-- Fairfax, VA, U.S.A.
-- =====================================================================

library ieee;
use ieee.std_logic_1164.all;

package sha3_hamsi_256cons is
	type gen256_type is array (0 to 15, 0 to 127) of std_logic_vector(1 downto 0);
	constant generator256 : gen256_type := (
	("01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", "01", "01", "11", "00", "00", "11", "11", "11", "11", "00", "00", "10", "00", "00",
	"11", "00", "10", "11", "10", "10", "01", "00", "10", "10", "11", "00", "11", "00", "00", "01", "00", "10", "01", "10", "11", "11", "11", "01", "10", "11", "11", "00", "01", "01", "01",
	"11", "01", "01", "01", "01", "00", "00", "11", "00", "00", "00", "11", "01", "11", "11", "10", "10", "10", "11", "00", "00", "10", "10", "11", "00", "01", "01", "10", "00", "01", "10",
	"01", "11", "00", "01", "10", "11", "01", "00", "01", "10", "01", "11", "11", "11", "11", "11", "10", "01", "01", "00", "10", "11", "10", "01", "00", "10", "11", "01", "01", "00", "10",
	"11", "11", "10", "00"),
	("00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "10", "11", "11", "00", "10", "01", "01", "01", "11", "00", "01", "10", "00",
	"10", "11", "01", "00", "10", "11", "01", "01", "01", "11", "00", "11", "10", "11", "00", "11", "01", "01", "01", "00", "00", "01", "01", "00", "00", "00", "01", "11", "11", "10", "10",
	"11", "00", "10", "10", "10", "01", "00", "10", "11", "00", "00", "10", "00", "11", "01", "10", "11", "11", "00", "11", "00", "01", "11", "00", "11", "11", "10", "00", "10", "11", "00",
	"01", "11", "11", "11", "00", "00", "00", "01", "11", "00", "01", "11", "01", "01", "01", "01", "10", "01", "10", "01", "01", "00", "10", "01", "01", "01", "00", "00", "10", "01", "01",
	"00", "01", "01", "10"),
	("00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "10", "10", "00", "11", "11", "10", "00", "11", "11", "01", "11", "01", "01", "10",
	"10", "10", "10", "11", "01", "11", "00", "01", "00", "00", "01", "00", "01", "10", "11", "11", "11", "00", "10", "00", "10", "10", "11", "10", "01", "10", "10", "01", "00", "00", "01",
	"00", "10", "11", "01", "01", "10", "01", "10", "10", "11", "00", "10", "01", "10", "01", "00", "11", "10", "01", "00", "11", "01", "00", "01", "00", "00", "00", "11", "00", "01", "10",
	"11", "11", "11", "00", "10", "10", "11", "00", "10", "10", "11", "11", "01", "11", "11", "11", "00", "01", "10", "10", "00", "11", "01", "01", "01", "00", "11", "11", "11", "10", "00",
	"11", "10", "00", "01"),
	("00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "10", "10", "00", "11", "11", "10", "00", "11", "11", "01", "11", "01", "01",
	"10", "10", "10", "10", "11", "01", "11", "00", "01", "00", "00", "01", "00", "01", "10", "11", "11", "11", "00", "10", "00", "10", "10", "11", "10", "01", "10", "10", "01", "00", "00",
	"01", "10", "10", "11", "01", "01", "10", "01", "10", "10", "11", "00", "10", "01", "10", "01", "00", "11", "10", "01", "00", "11", "01", "00", "01", "00", "00", "00", "11", "00", "01",
	"10", "11", "11", "11", "00", "10", "10", "11", "00", "10", "10", "11", "11", "01", "11", "11", "11", "00", "01", "10", "10", "00", "11", "01", "01", "01", "00", "11", "11", "11", "10",
	"00", "11", "01", "00"),
	("00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", "01", "00", "01", "10", "00", "00", "00", "01", "11", "11", "11", "11", "11", "01",
	"10", "10", "00", "01", "00", "01", "00", "11", "10", "11", "11", "00", "10", "00", "01", "11", "11", "01", "10", "10", "01", "11", "01", "11", "01", "01", "10", "10", "11", "00", "01",
	"11", "10", "11", "11", "10", "01", "01", "01", "01", "10", "10", "00", "01", "01", "10", "00", "11", "10", "00", "10", "01", "10", "01", "10", "00", "00", "01", "10", "00", "10", "10",
	"00", "01", "11", "10", "01", "11", "11", "10", "10", "10", "11", "01", "00", "00", "10", "00", "01", "10", "01", "01", "00", "01", "10", "10", "01", "11", "10", "01", "10", "11", "01",
	"01", "11", "11", "01"),
	("00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "01", "10", "10", "01", "10", "10", "10", "10", "11", "11", "11", "10", "11", "11",
	"11", "10", "11", "10", "00", "01", "10", "00", "10", "11", "01", "11", "10", "10", "00", "10", "11", "10", "10", "11", "00", "11", "01", "10", "10", "11", "11", "10", "01", "00", "11",
	"11", "00", "01", "00", "00", "10", "01", "11", "01", "01", "10", "00", "11", "11", "11", "11", "01", "10", "00", "00", "10", "00", "11", "11", "10", "11", "11", "00", "10", "11", "11",
	"01", "10", "01", "00", "11", "11", "00", "11", "01", "11", "01", "01", "11", "10", "10", "00", "01", "10", "01", "01", "00", "10", "00", "01", "10", "00", "01", "01", "10", "10", "10",
	"11", "11", "10", "11"),
	("00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "10", "10", "00", "10", "01", "00", "00", "00", "00", "11", "11", "10", "10", "11",
	"01", "11", "11", "01", "11", "01", "10", "10", "01", "11", "01", "01", "01", "10", "10", "11", "10", "10", "01", "11", "01", "10", "01", "10", "11", "00", "01", "11", "01", "10", "11",
	"01", "00", "11", "10", "11", "00", "10", "11", "11", "01", "01", "00", "11", "01", "01", "10", "10", "00", "00", "00", "00", "11", "01", "01", "11", "01", "00", "10", "00", "01", "10",
	"00", "11", "10", "10", "01", "01", "00", "00", "00", "00", "00", "11", "11", "01", "00", "00", "01", "10", "01", "01", "00", "10", "11", "11", "01", "11", "10", "10", "10", "10", "11",
	"00", "01", "10", "10"),
	("00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "10", "00", "11", "01", "00", "10", "10", "11", "11", "11", "00", "11", "01", "10", "10",
	"00", "01", "01", "00", "11", "01", "00", "10", "00", "11", "00", "01", "10", "01", "10", "11", "11", "00", "11", "11", "00", "10", "01", "00", "00", "00", "11", "01", "10", "00", "11",
	"00", "00", "01", "10", "11", "11", "00", "01", "11", "11", "01", "10", "01", "00", "10", "11", "00", "00", "11", "00", "00", "10", "01", "10", "01", "10", "00", "10", "10", "01", "11",
	"11", "11", "11", "11", "00", "10", "00", "00", "01", "10", "01", "11", "00", "00", "10", "11", "10", "00", "11", "01", "11", "11", "00", "10", "11", "11", "00", "11", "11", "10", "00",
	"00", "11", "00", "10"),
	("00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "00", "10", "00", "11", "01", "00", "10", "10", "11", "11", "11", "00", "11", "01", "10",
	"10", "00", "01", "01", "00", "11", "01", "00", "10", "00", "11", "00", "01", "10", "01", "10", "11", "11", "00", "11", "11", "00", "10", "01", "00", "00", "00", "11", "01", "10", "00",
	"11", "11", "00", "01", "10", "11", "11", "00", "01", "11", "11", "01", "10", "01", "00", "10", "11", "00", "00", "11", "00", "00", "10", "01", "10", "01", "10", "00", "10", "10", "01",
	"11", "11", "11", "11", "11", "00", "10", "00", "00", "01", "10", "01", "11", "00", "00", "10", "11", "10", "00", "11", "01", "11", "11", "00", "10", "11", "11", "00", "11", "11", "10",
	"00", "00", "11", "00"),
	("00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "00", "01", "11", "01", "10", "11", "01", "10", "00", "00", "01", "11", "11", "01", "11", "01",
	"00", "10", "01", "11", "00", "01", "00", "01", "01", "11", "10", "11", "10", "01", "10", "10", "10", "10", "00", "01", "01", "01", "10", "01", "00", "10", "10", "00", "00", "10", "01",
	"10", "11", "00", "11", "10", "10", "11", "01", "00", "01", "11", "01", "10", "00", "11", "01", "11", "10", "10", "00", "11", "01", "01", "00", "01", "01", "10", "11", "00", "01", "11",
	"10", "01", "11", "00", "10", "01", "11", "10", "11", "01", "10", "00", "11", "01", "10", "10", "11", "00", "01", "00", "10", "11", "10", "00", "00", "11", "01", "00", "11", "11", "10",
	"00", "10", "11", "11"),
	("00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "11", "11", "01", "00", "10", "11", "00", "11", "01", "01", "01", "11", "00", "01", "11",
	"00", "00", "01", "00", "00", "11", "11", "00", "10", "10", "10", "10", "10", "10", "01", "00", "10", "01", "00", "11", "00", "00", "00", "00", "10", "01", "11", "10", "10", "10", "00",
	"00", "00", "01", "10", "01", "10", "10", "10", "01", "00", "01", "10", "11", "11", "01", "00", "10", "00", "11", "10", "00", "00", "10", "00", "00", "11", "11", "01", "11", "10", "10",
	"01", "11", "01", "01", "11", "11", "11", "11", "00", "00", "11", "11", "01", "10", "00", "11", "01", "01", "10", "01", "11", "11", "00", "00", "00", "11", "10", "11", "10", "11", "00",
	"11", "01", "01", "11"),
	("00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "11", "11", "01", "00", "10", "11", "00", "11", "01", "01", "01", "11", "00", "01",
	"11", "00", "00", "01", "00", "00", "11", "11", "00", "10", "10", "10", "10", "10", "10", "01", "00", "10", "01", "00", "11", "00", "00", "00", "00", "10", "01", "11", "10", "10", "10",
	"00", "01", "00", "01", "10", "01", "10", "10", "10", "01", "00", "01", "10", "11", "11", "01", "00", "10", "00", "11", "10", "00", "00", "10", "00", "00", "11", "11", "01", "11", "10",
	"10", "01", "11", "01", "01", "11", "11", "11", "11", "00", "00", "11", "11", "01", "10", "00", "11", "01", "01", "10", "01", "11", "11", "00", "00", "00", "11", "10", "11", "10", "11",
	"00", "11", "01", "01"),
	("00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "00", "00", "00", "11", "11", "01", "00", "10", "11", "00", "11", "01", "01", "01", "11", "00",
	"01", "11", "00", "00", "01", "00", "00", "11", "11", "00", "10", "10", "10", "10", "10", "10", "01", "00", "10", "01", "00", "11", "00", "00", "00", "00", "10", "01", "11", "10", "10",
	"10", "11", "01", "00", "01", "10", "01", "10", "10", "10", "01", "00", "01", "10", "11", "11", "01", "00", "10", "00", "11", "10", "00", "00", "10", "00", "00", "11", "11", "01", "11",
	"10", "10", "01", "11", "01", "01", "11", "11", "11", "11", "00", "00", "11", "11", "01", "10", "00", "11", "01", "01", "10", "01", "11", "11", "00", "00", "00", "11", "10", "11", "10",
	"11", "00", "00", "01"),
	("00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "00", "11", "10", "10", "10", "11", "01", "01", "11", "10", "01", "11", "01", "10", "01", "11",
	"01", "01", "00", "01", "11", "10", "10", "00", "00", "00", "01", "10", "11", "10", "10", "00", "10", "10", "10", "01", "00", "01", "10", "10", "11", "01", "01", "10", "11", "01", "00",
	"11", "10", "01", "11", "10", "01", "10", "00", "10", "10", "10", "00", "10", "00", "11", "00", "00", "10", "01", "10", "00", "00", "01", "01", "00", "00", "10", "11", "11", "01", "10",
	"01", "11", "10", "11", "00", "00", "11", "11", "01", "00", "01", "01", "01", "10", "10", "00", "01", "10", "01", "01", "10", "11", "10", "01", "11", "11", "01", "10", "01", "10", "00",
	"11", "10", "01", "00"),
	("00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "00", "01", "00", "01", "00", "10", "11", "11", "11", "01", "00", "01", "11", "00", "10", "01",
	"01", "01", "00", "10", "00", "10", "01", "10", "01", "01", "10", "01", "00", "11", "10", "01", "00", "11", "01", "11", "11", "10", "11", "01", "11", "01", "11", "01", "01", "00", "10",
	"10", "01", "01", "10", "00", "10", "01", "00", "00", "10", "10", "00", "11", "00", "10", "10", "01", "01", "00", "01", "10", "01", "01", "11", "01", "11", "11", "11", "11", "00", "00",
	"01", "11", "11", "01", "10", "10", "11", "11", "00", "00", "11", "11", "11", "11", "00", "00", "01", "10", "01", "01", "00", "00", "10", "01", "01", "10", "01", "10", "01", "01", "11",
	"10", "01", "00", "01"),
	("00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", "11", "11", "10", "00", "00", "10", "10", "10", "10", "00", "00", "01", "00", "00", "10",
	"00", "01", "10", "01", "01", "11", "00", "01", "01", "10", "00", "10", "00", "00", "11", "00", "01", "11", "01", "10", "10", "10", "11", "01", "10", "10", "00", "11", "11", "11", "10",
	"11", "11", "11", "11", "00", "00", "10", "00", "00", "00", "10", "11", "10", "10", "01", "01", "01", "10", "00", "00", "01", "01", "10", "00", "11", "11", "01", "00", "11", "01", "11",
	"10", "00", "11", "01", "10", "11", "00", "11", "01", "11", "10", "10", "10", "10", "10", "01", "11", "11", "00", "01", "10", "01", "11", "00", "01", "10", "11", "11", "00", "01", "10",
	"10", "11", "00", "00"));
	
	TYPE vec_array IS ARRAY (0 to 255, 0 to 7) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	TYPE vector_array IS ARRAY (0 to 3) OF vec_array;
-- constans used in P
	CONSTANT g256 : vector_array := (
	(
		(x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000"), 
		(x"74951000", x"5A2B467E", x"88FD1D2B", x"1EE68292", x"CBA90000", x"90273769", x"BBDCF407", x"D0F4AF61"), 
		(x"CBA90000", x"90273769", x"BBDCF407", x"D0F4AF61", x"BF3C1000", x"CA0C7117", x"3321E92C", x"CE122DF3"), 
		(x"BF3C1000", x"CA0C7117", x"3321E92C", x"CE122DF3", x"74951000", x"5A2B467E", x"88FD1D2B", x"1EE68292"), 
		(x"E92A2000", x"B4578CFC", x"11FA3A57", x"3DC90524", x"97530000", x"204F6ED3", x"77B9E80F", x"A1EC5EC1"), 
		(x"9DBF3000", x"EE7CCA82", x"9907277C", x"232F87B6", x"5CFA0000", x"B06859BA", x"CC651C08", x"7118F1A0"), 
		(x"22832000", x"2470BB95", x"AA26CE50", x"ED3DAA45", x"286F1000", x"EA431FC4", x"44980123", x"6FFE7332"), 
		(x"56163000", x"7E5BFDEB", x"22DBD37B", x"F3DB28D7", x"E3C61000", x"7A6428AD", x"FF44F524", x"BF0ADC53"), 
		(x"97530000", x"204F6ED3", x"77B9E80F", x"A1EC5EC1", x"7E792000", x"9418E22F", x"6643D258", x"9C255BE5"), 
		(x"E3C61000", x"7A6428AD", x"FF44F524", x"BF0ADC53", x"B5D02000", x"043FD546", x"DD9F265F", x"4CD1F484"), 
		(x"5CFA0000", x"B06859BA", x"CC651C08", x"7118F1A0", x"C1453000", x"5E149338", x"55623B74", x"52377616"), 
		(x"286F1000", x"EA431FC4", x"44980123", x"6FFE7332", x"0AEC3000", x"CE33A451", x"EEBECF73", x"82C3D977"), 
		(x"7E792000", x"9418E22F", x"6643D258", x"9C255BE5", x"E92A2000", x"B4578CFC", x"11FA3A57", x"3DC90524"), 
		(x"0AEC3000", x"CE33A451", x"EEBECF73", x"82C3D977", x"22832000", x"2470BB95", x"AA26CE50", x"ED3DAA45"), 
		(x"B5D02000", x"043FD546", x"DD9F265F", x"4CD1F484", x"56163000", x"7E5BFDEB", x"22DBD37B", x"F3DB28D7"), 
		(x"C1453000", x"5E149338", x"55623B74", x"52377616", x"9DBF3000", x"EE7CCA82", x"9907277C", x"232F87B6"), 
		(x"121B4000", x"5B17D9E8", x"8DFACFAB", x"CE36CC72", x"E6570000", x"4BB33A25", x"848598BA", x"1041003E"), 
		(x"668E5000", x"013C9F96", x"0507D280", x"D0D04EE0", x"2DFE0000", x"DB940D4C", x"3F596CBD", x"C0B5AF5F"), 
		(x"D9B24000", x"CB30EE81", x"36263BAC", x"1EC26313", x"596B1000", x"81BF4B32", x"B7A47196", x"DE532DCD"), 
		(x"AD275000", x"911BA8FF", x"BEDB2687", x"0024E181", x"92C21000", x"11987C5B", x"0C788591", x"0EA782AC"), 
		(x"FB316000", x"EF405514", x"9C00F5FC", x"F3FFC956", x"71040000", x"6BFC54F6", x"F33C70B5", x"B1AD5EFF"), 
		(x"8FA47000", x"B56B136A", x"14FDE8D7", x"ED194BC4", x"BAAD0000", x"FBDB639F", x"48E084B2", x"6159F19E"), 
		(x"30986000", x"7F67627D", x"27DC01FB", x"230B6637", x"CE381000", x"A1F025E1", x"C01D9999", x"7FBF730C"), 
		(x"440D7000", x"254C2403", x"AF211CD0", x"3DEDE4A5", x"05911000", x"31D71288", x"7BC16D9E", x"AF4BDC6D"), 
		(x"85484000", x"7B58B73B", x"FA4327A4", x"6FDA92B3", x"982E2000", x"DFABD80A", x"E2C64AE2", x"8C645BDB"), 
		(x"F1DD5000", x"2173F145", x"72BE3A8F", x"713C1021", x"53872000", x"4F8CEF63", x"591ABEE5", x"5C90F4BA"), 
		(x"4EE14000", x"EB7F8052", x"419FD3A3", x"BF2E3DD2", x"27123000", x"15A7A91D", x"D1E7A3CE", x"42767628"), 
		(x"3A745000", x"B154C62C", x"C962CE88", x"A1C8BF40", x"ECBB3000", x"85809E74", x"6A3B57C9", x"9282D949"), 
		(x"6C626000", x"CF0F3BC7", x"EBB91DF3", x"52139797", x"0F7D2000", x"FFE4B6D9", x"957FA2ED", x"2D88051A"), 
		(x"18F77000", x"95247DB9", x"634400D8", x"4CF51505", x"C4D42000", x"6FC381B0", x"2EA356EA", x"FD7CAA7B"), 
		(x"A7CB6000", x"5F280CAE", x"5065E9F4", x"82E738F6", x"B0413000", x"35E8C7CE", x"A65E4BC1", x"E39A28E9"), 
		(x"D35E7000", x"05034AD0", x"D898F4DF", x"9C01BA64", x"7BE83000", x"A5CFF0A7", x"1D82BFC6", x"336E8788"), 
		(x"E6570000", x"4BB33A25", x"848598BA", x"1041003E", x"F44C4000", x"10A4E3CD", x"097F5711", x"DE77CC4C"), 
		(x"92C21000", x"11987C5B", x"0C788591", x"0EA782AC", x"3FE54000", x"8083D4A4", x"B2A3A316", x"0E83632D"), 
		(x"2DFE0000", x"DB940D4C", x"3F596CBD", x"C0B5AF5F", x"4B705000", x"DAA892DA", x"3A5EBE3D", x"1065E1BF"), 
		(x"596B1000", x"81BF4B32", x"B7A47196", x"DE532DCD", x"80D95000", x"4A8FA5B3", x"81824A3A", x"C0914EDE"), 
		(x"0F7D2000", x"FFE4B6D9", x"957FA2ED", x"2D88051A", x"631F4000", x"30EB8D1E", x"7EC6BF1E", x"7F9B928D"), 
		(x"7BE83000", x"A5CFF0A7", x"1D82BFC6", x"336E8788", x"A8B64000", x"A0CCBA77", x"C51A4B19", x"AF6F3DEC"), 
		(x"C4D42000", x"6FC381B0", x"2EA356EA", x"FD7CAA7B", x"DC235000", x"FAE7FC09", x"4DE75632", x"B189BF7E"), 
		(x"B0413000", x"35E8C7CE", x"A65E4BC1", x"E39A28E9", x"178A5000", x"6AC0CB60", x"F63BA235", x"617D101F"), 
		(x"71040000", x"6BFC54F6", x"F33C70B5", x"B1AD5EFF", x"8A356000", x"84BC01E2", x"6F3C8549", x"425297A9"), 
		(x"05911000", x"31D71288", x"7BC16D9E", x"AF4BDC6D", x"419C6000", x"149B368B", x"D4E0714E", x"92A638C8"), 
		(x"BAAD0000", x"FBDB639F", x"48E084B2", x"6159F19E", x"35097000", x"4EB070F5", x"5C1D6C65", x"8C40BA5A"), 
		(x"CE381000", x"A1F025E1", x"C01D9999", x"7FBF730C", x"FEA07000", x"DE97479C", x"E7C19862", x"5CB4153B"), 
		(x"982E2000", x"DFABD80A", x"E2C64AE2", x"8C645BDB", x"1D666000", x"A4F36F31", x"18856D46", x"E3BEC968"), 
		(x"ECBB3000", x"85809E74", x"6A3B57C9", x"9282D949", x"D6CF6000", x"34D45858", x"A3599941", x"334A6609"), 
		(x"53872000", x"4F8CEF63", x"591ABEE5", x"5C90F4BA", x"A25A7000", x"6EFF1E26", x"2BA4846A", x"2DACE49B"), 
		(x"27123000", x"15A7A91D", x"D1E7A3CE", x"42767628", x"69F37000", x"FED8294F", x"9078706D", x"FD584BFA"), 
		(x"F44C4000", x"10A4E3CD", x"097F5711", x"DE77CC4C", x"121B4000", x"5B17D9E8", x"8DFACFAB", x"CE36CC72"), 
		(x"80D95000", x"4A8FA5B3", x"81824A3A", x"C0914EDE", x"D9B24000", x"CB30EE81", x"36263BAC", x"1EC26313"), 
		(x"3FE54000", x"8083D4A4", x"B2A3A316", x"0E83632D", x"AD275000", x"911BA8FF", x"BEDB2687", x"0024E181"), 
		(x"4B705000", x"DAA892DA", x"3A5EBE3D", x"1065E1BF", x"668E5000", x"013C9F96", x"0507D280", x"D0D04EE0"), 
		(x"1D666000", x"A4F36F31", x"18856D46", x"E3BEC968", x"85484000", x"7B58B73B", x"FA4327A4", x"6FDA92B3"), 
		(x"69F37000", x"FED8294F", x"9078706D", x"FD584BFA", x"4EE14000", x"EB7F8052", x"419FD3A3", x"BF2E3DD2"), 
		(x"D6CF6000", x"34D45858", x"A3599941", x"334A6609", x"3A745000", x"B154C62C", x"C962CE88", x"A1C8BF40"), 
		(x"A25A7000", x"6EFF1E26", x"2BA4846A", x"2DACE49B", x"F1DD5000", x"2173F145", x"72BE3A8F", x"713C1021"), 
		(x"631F4000", x"30EB8D1E", x"7EC6BF1E", x"7F9B928D", x"6C626000", x"CF0F3BC7", x"EBB91DF3", x"52139797"), 
		(x"178A5000", x"6AC0CB60", x"F63BA235", x"617D101F", x"A7CB6000", x"5F280CAE", x"5065E9F4", x"82E738F6"), 
		(x"A8B64000", x"A0CCBA77", x"C51A4B19", x"AF6F3DEC", x"D35E7000", x"05034AD0", x"D898F4DF", x"9C01BA64"), 
		(x"DC235000", x"FAE7FC09", x"4DE75632", x"B189BF7E", x"18F77000", x"95247DB9", x"634400D8", x"4CF51505"), 
		(x"8A356000", x"84BC01E2", x"6F3C8549", x"425297A9", x"FB316000", x"EF405514", x"9C00F5FC", x"F3FFC956"), 
		(x"FEA07000", x"DE97479C", x"E7C19862", x"5CB4153B", x"30986000", x"7F67627D", x"27DC01FB", x"230B6637"), 
		(x"419C6000", x"149B368B", x"D4E0714E", x"92A638C8", x"440D7000", x"254C2403", x"AF211CD0", x"3DEDE4A5"), 
		(x"35097000", x"4EB070F5", x"5C1D6C65", x"8C40BA5A", x"8FA47000", x"B56B136A", x"14FDE8D7", x"ED194BC4"), 
		(x"E4788000", x"859673C1", x"B5FB2452", x"29CC5EDF", x"045F0000", x"9C4A93C9", x"62FC79D0", x"731EBDC2"), 
		(x"90ED9000", x"DFBD35BF", x"3D063979", x"372ADC4D", x"CFF60000", x"0C6DA4A0", x"D9208DD7", x"A3EA12A3"), 
		(x"2FD18000", x"15B144A8", x"0E27D055", x"F938F1BE", x"BB631000", x"5646E2DE", x"51DD90FC", x"BD0C9031"), 
		(x"5B449000", x"4F9A02D6", x"86DACD7E", x"E7DE732C", x"70CA1000", x"C661D5B7", x"EA0164FB", x"6DF83F50"), 
		(x"0D52A000", x"31C1FF3D", x"A4011E05", x"14055BFB", x"930C0000", x"BC05FD1A", x"154591DF", x"D2F2E303"), 
		(x"79C7B000", x"6BEAB943", x"2CFC032E", x"0AE3D969", x"58A50000", x"2C22CA73", x"AE9965D8", x"02064C62"), 
		(x"C6FBA000", x"A1E6C854", x"1FDDEA02", x"C4F1F49A", x"2C301000", x"76098C0D", x"266478F3", x"1CE0CEF0"), 
		(x"B26EB000", x"FBCD8E2A", x"9720F729", x"DA177608", x"E7991000", x"E62EBB64", x"9DB88CF4", x"CC146191"), 
		(x"732B8000", x"A5D91D12", x"C242CC5D", x"8820001E", x"7A262000", x"085271E6", x"04BFAB88", x"EF3BE627"), 
		(x"07BE9000", x"FFF25B6C", x"4ABFD176", x"96C6828C", x"B18F2000", x"9875468F", x"BF635F8F", x"3FCF4946"), 
		(x"B8828000", x"35FE2A7B", x"799E385A", x"58D4AF7F", x"C51A3000", x"C25E00F1", x"379E42A4", x"2129CBD4"), 
		(x"CC179000", x"6FD56C05", x"F1632571", x"46322DED", x"0EB33000", x"52793798", x"8C42B6A3", x"F1DD64B5"), 
		(x"9A01A000", x"118E91EE", x"D3B8F60A", x"B5E9053A", x"ED752000", x"281D1F35", x"73064387", x"4ED7B8E6"), 
		(x"EE94B000", x"4BA5D790", x"5B45EB21", x"AB0F87A8", x"26DC2000", x"B83A285C", x"C8DAB780", x"9E231787"), 
		(x"51A8A000", x"81A9A687", x"6864020D", x"651DAA5B", x"52493000", x"E2116E22", x"4027AAAB", x"80C59515"), 
		(x"253DB000", x"DB82E0F9", x"E0991F26", x"7BFB28C9", x"99E03000", x"7236594B", x"FBFB5EAC", x"50313A74"), 
		(x"F663C000", x"DE81AA29", x"3801EBF9", x"E7FA92AD", x"E2080000", x"D7F9A9EC", x"E679E16A", x"635FBDFC"), 
		(x"82F6D000", x"84AAEC57", x"B0FCF6D2", x"F91C103F", x"29A10000", x"47DE9E85", x"5DA5156D", x"B3AB129D"), 
		(x"3DCAC000", x"4EA69D40", x"83DD1FFE", x"370E3DCC", x"5D341000", x"1DF5D8FB", x"D5580846", x"AD4D900F"), 
		(x"495FD000", x"148DDB3E", x"0B2002D5", x"29E8BF5E", x"969D1000", x"8DD2EF92", x"6E84FC41", x"7DB93F6E"), 
		(x"1F49E000", x"6AD626D5", x"29FBD1AE", x"DA339789", x"755B0000", x"F7B6C73F", x"91C00965", x"C2B3E33D"), 
		(x"6BDCF000", x"30FD60AB", x"A106CC85", x"C4D5151B", x"BEF20000", x"6791F056", x"2A1CFD62", x"12474C5C"), 
		(x"D4E0E000", x"FAF111BC", x"922725A9", x"0AC738E8", x"CA671000", x"3DBAB628", x"A2E1E049", x"0CA1CECE"), 
		(x"A075F000", x"A0DA57C2", x"1ADA3882", x"1421BA7A", x"01CE1000", x"AD9D8141", x"193D144E", x"DC5561AF"), 
		(x"6130C000", x"FECEC4FA", x"4FB803F6", x"4616CC6C", x"9C712000", x"43E14BC3", x"803A3332", x"FF7AE619"), 
		(x"15A5D000", x"A4E58284", x"C7451EDD", x"58F04EFE", x"57D82000", x"D3C67CAA", x"3BE6C735", x"2F8E4978"), 
		(x"AA99C000", x"6EE9F393", x"F464F7F1", x"96E2630D", x"234D3000", x"89ED3AD4", x"B31BDA1E", x"3168CBEA"), 
		(x"DE0CD000", x"34C2B5ED", x"7C99EADA", x"8804E19F", x"E8E43000", x"19CA0DBD", x"08C72E19", x"E19C648B"), 
		(x"881AE000", x"4A994806", x"5E4239A1", x"7BDFC948", x"0B222000", x"63AE2510", x"F783DB3D", x"5E96B8D8"), 
		(x"FC8FF000", x"10B20E78", x"D6BF248A", x"65394BDA", x"C08B2000", x"F3891279", x"4C5F2F3A", x"8E6217B9"), 
		(x"43B3E000", x"DABE7F6F", x"E59ECDA6", x"AB2B6629", x"B41E3000", x"A9A25407", x"C4A23211", x"9084952B"), 
		(x"3726F000", x"80953911", x"6D63D08D", x"B5CDE4BB", x"7FB73000", x"3985636E", x"7F7EC616", x"40703A4A"), 
		(x"022F8000", x"CE2549E4", x"317EBCE8", x"398D5EE1", x"F0134000", x"8CEE7004", x"6B832EC1", x"AD69718E"), 
		(x"76BA9000", x"940E0F9A", x"B983A1C3", x"276BDC73", x"3BBA4000", x"1CC9476D", x"D05FDAC6", x"7D9DDEEF"), 
		(x"C9868000", x"5E027E8D", x"8AA248EF", x"E979F180", x"4F2F5000", x"46E20113", x"58A2C7ED", x"637B5C7D"), 
		(x"BD139000", x"042938F3", x"025F55C4", x"F79F7312", x"84865000", x"D6C5367A", x"E37E33EA", x"B38FF31C"), 
		(x"EB05A000", x"7A72C518", x"208486BF", x"04445BC5", x"67404000", x"ACA11ED7", x"1C3AC6CE", x"0C852F4F"), 
		(x"9F90B000", x"20598366", x"A8799B94", x"1AA2D957", x"ACE94000", x"3C8629BE", x"A7E632C9", x"DC71802E"), 
		(x"20ACA000", x"EA55F271", x"9B5872B8", x"D4B0F4A4", x"D87C5000", x"66AD6FC0", x"2F1B2FE2", x"C29702BC"), 
		(x"5439B000", x"B07EB40F", x"13A56F93", x"CA567636", x"13D55000", x"F68A58A9", x"94C7DBE5", x"1263ADDD"), 
		(x"957C8000", x"EE6A2737", x"46C754E7", x"98610020", x"8E6A6000", x"18F6922B", x"0DC0FC99", x"314C2A6B"), 
		(x"E1E99000", x"B4416149", x"CE3A49CC", x"868782B2", x"45C36000", x"88D1A542", x"B61C089E", x"E1B8850A"), 
		(x"5ED58000", x"7E4D105E", x"FD1BA0E0", x"4895AF41", x"31567000", x"D2FAE33C", x"3EE115B5", x"FF5E0798"), 
		(x"2A409000", x"24665620", x"75E6BDCB", x"56732DD3", x"FAFF7000", x"42DDD455", x"853DE1B2", x"2FAAA8F9"), 
		(x"7C56A000", x"5A3DABCB", x"573D6EB0", x"A5A80504", x"19396000", x"38B9FCF8", x"7A791496", x"90A074AA"), 
		(x"08C3B000", x"0016EDB5", x"DFC0739B", x"BB4E8796", x"D2906000", x"A89ECB91", x"C1A5E091", x"4054DBCB"), 
		(x"B7FFA000", x"CA1A9CA2", x"ECE19AB7", x"755CAA65", x"A6057000", x"F2B58DEF", x"4958FDBA", x"5EB25959"), 
		(x"C36AB000", x"9031DADC", x"641C879C", x"6BBA28F7", x"6DAC7000", x"6292BA86", x"F28409BD", x"8E46F638"), 
		(x"1034C000", x"9532900C", x"BC847343", x"F7BB9293", x"16444000", x"C75D4A21", x"EF06B67B", x"BD2871B0"), 
		(x"64A1D000", x"CF19D672", x"34796E68", x"E95D1001", x"DDED4000", x"577A7D48", x"54DA427C", x"6DDCDED1"), 
		(x"DB9DC000", x"0515A765", x"07588744", x"274F3DF2", x"A9785000", x"0D513B36", x"DC275F57", x"733A5C43"), 
		(x"AF08D000", x"5F3EE11B", x"8FA59A6F", x"39A9BF60", x"62D15000", x"9D760C5F", x"67FBAB50", x"A3CEF322"), 
		(x"F91EE000", x"21651CF0", x"AD7E4914", x"CA7297B7", x"81174000", x"E71224F2", x"98BF5E74", x"1CC42F71"), 
		(x"8D8BF000", x"7B4E5A8E", x"2583543F", x"D4941525", x"4ABE4000", x"7735139B", x"2363AA73", x"CC308010"), 
		(x"32B7E000", x"B1422B99", x"16A2BD13", x"1A8638D6", x"3E2B5000", x"2D1E55E5", x"AB9EB758", x"D2D60282"), 
		(x"4622F000", x"EB696DE7", x"9E5FA038", x"0460BA44", x"F5825000", x"BD39628C", x"1042435F", x"0222ADE3"), 
		(x"8767C000", x"B57DFEDF", x"CB3D9B4C", x"5657CC52", x"683D6000", x"5345A80E", x"89456423", x"210D2A55"), 
		(x"F3F2D000", x"EF56B8A1", x"43C08667", x"48B14EC0", x"A3946000", x"C3629F67", x"32999024", x"F1F98534"), 
		(x"4CCEC000", x"255AC9B6", x"70E16F4B", x"86A36333", x"D7017000", x"9949D919", x"BA648D0F", x"EF1F07A6"), 
		(x"385BD000", x"7F718FC8", x"F81C7260", x"9845E1A1", x"1CA87000", x"096EEE70", x"01B87908", x"3FEBA8C7"), 
		(x"6E4DE000", x"012A7223", x"DAC7A11B", x"6B9EC976", x"FF6E6000", x"730AC6DD", x"FEFC8C2C", x"80E17494"), 
		(x"1AD8F000", x"5B01345D", x"523ABC30", x"75784BE4", x"34C76000", x"E32DF1B4", x"4520782B", x"5015DBF5"), 
		(x"A5E4E000", x"910D454A", x"611B551C", x"BB6A6617", x"40527000", x"B906B7CA", x"CDDD6500", x"4EF35967"), 
		(x"D171F000", x"CB260334", x"E9E64837", x"A58CE485", x"8BFB7000", x"292180A3", x"76019107", x"9E07F606"), 
		(x"045F0000", x"9C4A93C9", x"62FC79D0", x"731EBDC2", x"E0278000", x"19DCE008", x"D7075D82", x"5AD2E31D"), 
		(x"70CA1000", x"C661D5B7", x"EA0164FB", x"6DF83F50", x"2B8E8000", x"89FBD761", x"6CDBA985", x"8A264C7C"), 
		(x"CFF60000", x"0C6DA4A0", x"D9208DD7", x"A3EA12A3", x"5F1B9000", x"D3D0911F", x"E426B4AE", x"94C0CEEE"), 
		(x"BB631000", x"5646E2DE", x"51DD90FC", x"BD0C9031", x"94B29000", x"43F7A676", x"5FFA40A9", x"4434618F"), 
		(x"ED752000", x"281D1F35", x"73064387", x"4ED7B8E6", x"77748000", x"39938EDB", x"A0BEB58D", x"FB3EBDDC"), 
		(x"99E03000", x"7236594B", x"FBFB5EAC", x"50313A74", x"BCDD8000", x"A9B4B9B2", x"1B62418A", x"2BCA12BD"), 
		(x"26DC2000", x"B83A285C", x"C8DAB780", x"9E231787", x"C8489000", x"F39FFFCC", x"939F5CA1", x"352C902F"), 
		(x"52493000", x"E2116E22", x"4027AAAB", x"80C59515", x"03E19000", x"63B8C8A5", x"2843A8A6", x"E5D83F4E"), 
		(x"930C0000", x"BC05FD1A", x"154591DF", x"D2F2E303", x"9E5EA000", x"8DC40227", x"B1448FDA", x"C6F7B8F8"), 
		(x"E7991000", x"E62EBB64", x"9DB88CF4", x"CC146191", x"55F7A000", x"1DE3354E", x"0A987BDD", x"16031799"), 
		(x"58A50000", x"2C22CA73", x"AE9965D8", x"02064C62", x"2162B000", x"47C87330", x"826566F6", x"08E5950B"), 
		(x"2C301000", x"76098C0D", x"266478F3", x"1CE0CEF0", x"EACBB000", x"D7EF4459", x"39B992F1", x"D8113A6A"), 
		(x"7A262000", x"085271E6", x"04BFAB88", x"EF3BE627", x"090DA000", x"AD8B6CF4", x"C6FD67D5", x"671BE639"), 
		(x"0EB33000", x"52793798", x"8C42B6A3", x"F1DD64B5", x"C2A4A000", x"3DAC5B9D", x"7D2193D2", x"B7EF4958"), 
		(x"B18F2000", x"9875468F", x"BF635F8F", x"3FCF4946", x"B631B000", x"67871DE3", x"F5DC8EF9", x"A909CBCA"), 
		(x"C51A3000", x"C25E00F1", x"379E42A4", x"2129CBD4", x"7D98B000", x"F7A02A8A", x"4E007AFE", x"79FD64AB"), 
		(x"16444000", x"C75D4A21", x"EF06B67B", x"BD2871B0", x"06708000", x"526FDA2D", x"5382C538", x"4A93E323"), 
		(x"62D15000", x"9D760C5F", x"67FBAB50", x"A3CEF322", x"CDD98000", x"C248ED44", x"E85E313F", x"9A674C42"), 
		(x"DDED4000", x"577A7D48", x"54DA427C", x"6DDCDED1", x"B94C9000", x"9863AB3A", x"60A32C14", x"8481CED0"), 
		(x"A9785000", x"0D513B36", x"DC275F57", x"733A5C43", x"72E59000", x"08449C53", x"DB7FD813", x"547561B1"), 
		(x"FF6E6000", x"730AC6DD", x"FEFC8C2C", x"80E17494", x"91238000", x"7220B4FE", x"243B2D37", x"EB7FBDE2"), 
		(x"8BFB7000", x"292180A3", x"76019107", x"9E07F606", x"5A8A8000", x"E2078397", x"9FE7D930", x"3B8B1283"), 
		(x"34C76000", x"E32DF1B4", x"4520782B", x"5015DBF5", x"2E1F9000", x"B82CC5E9", x"171AC41B", x"256D9011"), 
		(x"40527000", x"B906B7CA", x"CDDD6500", x"4EF35967", x"E5B69000", x"280BF280", x"ACC6301C", x"F5993F70"), 
		(x"81174000", x"E71224F2", x"98BF5E74", x"1CC42F71", x"7809A000", x"C6773802", x"35C11760", x"D6B6B8C6"), 
		(x"F5825000", x"BD39628C", x"1042435F", x"0222ADE3", x"B3A0A000", x"56500F6B", x"8E1DE367", x"064217A7"), 
		(x"4ABE4000", x"7735139B", x"2363AA73", x"CC308010", x"C735B000", x"0C7B4915", x"06E0FE4C", x"18A49535"), 
		(x"3E2B5000", x"2D1E55E5", x"AB9EB758", x"D2D60282", x"0C9CB000", x"9C5C7E7C", x"BD3C0A4B", x"C8503A54"), 
		(x"683D6000", x"5345A80E", x"89456423", x"210D2A55", x"EF5AA000", x"E63856D1", x"4278FF6F", x"775AE607"), 
		(x"1CA87000", x"096EEE70", x"01B87908", x"3FEBA8C7", x"24F3A000", x"761F61B8", x"F9A40B68", x"A7AE4966"), 
		(x"A3946000", x"C3629F67", x"32999024", x"F1F98534", x"5066B000", x"2C3427C6", x"71591643", x"B948CBF4"), 
		(x"D7017000", x"9949D919", x"BA648D0F", x"EF1F07A6", x"9BCFB000", x"BC1310AF", x"CA85E244", x"69BC6495"), 
		(x"E2080000", x"D7F9A9EC", x"E679E16A", x"635FBDFC", x"146BC000", x"097803C5", x"DE780A93", x"84A52F51"), 
		(x"969D1000", x"8DD2EF92", x"6E84FC41", x"7DB93F6E", x"DFC2C000", x"995F34AC", x"65A4FE94", x"54518030"), 
		(x"29A10000", x"47DE9E85", x"5DA5156D", x"B3AB129D", x"AB57D000", x"C37472D2", x"ED59E3BF", x"4AB702A2"), 
		(x"5D341000", x"1DF5D8FB", x"D5580846", x"AD4D900F", x"60FED000", x"535345BB", x"568517B8", x"9A43ADC3"), 
		(x"0B222000", x"63AE2510", x"F783DB3D", x"5E96B8D8", x"8338C000", x"29376D16", x"A9C1E29C", x"25497190"), 
		(x"7FB73000", x"3985636E", x"7F7EC616", x"40703A4A", x"4891C000", x"B9105A7F", x"121D169B", x"F5BDDEF1"), 
		(x"C08B2000", x"F3891279", x"4C5F2F3A", x"8E6217B9", x"3C04D000", x"E33B1C01", x"9AE00BB0", x"EB5B5C63"), 
		(x"B41E3000", x"A9A25407", x"C4A23211", x"9084952B", x"F7ADD000", x"731C2B68", x"213CFFB7", x"3BAFF302"), 
		(x"755B0000", x"F7B6C73F", x"91C00965", x"C2B3E33D", x"6A12E000", x"9D60E1EA", x"B83BD8CB", x"188074B4"), 
		(x"01CE1000", x"AD9D8141", x"193D144E", x"DC5561AF", x"A1BBE000", x"0D47D683", x"03E72CCC", x"C874DBD5"), 
		(x"BEF20000", x"6791F056", x"2A1CFD62", x"12474C5C", x"D52EF000", x"576C90FD", x"8B1A31E7", x"D6925947"), 
		(x"CA671000", x"3DBAB628", x"A2E1E049", x"0CA1CECE", x"1E87F000", x"C74BA794", x"30C6C5E0", x"0666F626"), 
		(x"9C712000", x"43E14BC3", x"803A3332", x"FF7AE619", x"FD41E000", x"BD2F8F39", x"CF8230C4", x"B96C2A75"), 
		(x"E8E43000", x"19CA0DBD", x"08C72E19", x"E19C648B", x"36E8E000", x"2D08B850", x"745EC4C3", x"69988514"), 
		(x"57D82000", x"D3C67CAA", x"3BE6C735", x"2F8E4978", x"427DF000", x"7723FE2E", x"FCA3D9E8", x"777E0786"), 
		(x"234D3000", x"89ED3AD4", x"B31BDA1E", x"3168CBEA", x"89D4F000", x"E704C947", x"477F2DEF", x"A78AA8E7"), 
		(x"F0134000", x"8CEE7004", x"6B832EC1", x"AD69718E", x"F23CC000", x"42CB39E0", x"5AFD9229", x"94E42F6F"), 
		(x"84865000", x"D6C5367A", x"E37E33EA", x"B38FF31C", x"3995C000", x"D2EC0E89", x"E121662E", x"4410800E"), 
		(x"3BBA4000", x"1CC9476D", x"D05FDAC6", x"7D9DDEEF", x"4D00D000", x"88C748F7", x"69DC7B05", x"5AF6029C"), 
		(x"4F2F5000", x"46E20113", x"58A2C7ED", x"637B5C7D", x"86A9D000", x"18E07F9E", x"D2008F02", x"8A02ADFD"), 
		(x"19396000", x"38B9FCF8", x"7A791496", x"90A074AA", x"656FC000", x"62845733", x"2D447A26", x"350871AE"), 
		(x"6DAC7000", x"6292BA86", x"F28409BD", x"8E46F638", x"AEC6C000", x"F2A3605A", x"96988E21", x"E5FCDECF"), 
		(x"D2906000", x"A89ECB91", x"C1A5E091", x"4054DBCB", x"DA53D000", x"A8882624", x"1E65930A", x"FB1A5C5D"), 
		(x"A6057000", x"F2B58DEF", x"4958FDBA", x"5EB25959", x"11FAD000", x"38AF114D", x"A5B9670D", x"2BEEF33C"), 
		(x"67404000", x"ACA11ED7", x"1C3AC6CE", x"0C852F4F", x"8C45E000", x"D6D3DBCF", x"3CBE4071", x"08C1748A"), 
		(x"13D55000", x"F68A58A9", x"94C7DBE5", x"1263ADDD", x"47ECE000", x"46F4ECA6", x"8762B476", x"D835DBEB"), 
		(x"ACE94000", x"3C8629BE", x"A7E632C9", x"DC71802E", x"3379F000", x"1CDFAAD8", x"0F9FA95D", x"C6D35979"), 
		(x"D87C5000", x"66AD6FC0", x"2F1B2FE2", x"C29702BC", x"F8D0F000", x"8CF89DB1", x"B4435D5A", x"1627F618"), 
		(x"8E6A6000", x"18F6922B", x"0DC0FC99", x"314C2A6B", x"1B16E000", x"F69CB51C", x"4B07A87E", x"A92D2A4B"), 
		(x"FAFF7000", x"42DDD455", x"853DE1B2", x"2FAAA8F9", x"D0BFE000", x"66BB8275", x"F0DB5C79", x"79D9852A"), 
		(x"45C36000", x"88D1A542", x"B61C089E", x"E1B8850A", x"A42AF000", x"3C90C40B", x"78264152", x"673F07B8"), 
		(x"31567000", x"D2FAE33C", x"3EE115B5", x"FF5E0798", x"6F83F000", x"ACB7F362", x"C3FAB555", x"B7CBA8D9"), 
		(x"E0278000", x"19DCE008", x"D7075D82", x"5AD2E31D", x"E4788000", x"859673C1", x"B5FB2452", x"29CC5EDF"), 
		(x"94B29000", x"43F7A676", x"5FFA40A9", x"4434618F", x"2FD18000", x"15B144A8", x"0E27D055", x"F938F1BE"), 
		(x"2B8E8000", x"89FBD761", x"6CDBA985", x"8A264C7C", x"5B449000", x"4F9A02D6", x"86DACD7E", x"E7DE732C"), 
		(x"5F1B9000", x"D3D0911F", x"E426B4AE", x"94C0CEEE", x"90ED9000", x"DFBD35BF", x"3D063979", x"372ADC4D"), 
		(x"090DA000", x"AD8B6CF4", x"C6FD67D5", x"671BE639", x"732B8000", x"A5D91D12", x"C242CC5D", x"8820001E"), 
		(x"7D98B000", x"F7A02A8A", x"4E007AFE", x"79FD64AB", x"B8828000", x"35FE2A7B", x"799E385A", x"58D4AF7F"), 
		(x"C2A4A000", x"3DAC5B9D", x"7D2193D2", x"B7EF4958", x"CC179000", x"6FD56C05", x"F1632571", x"46322DED"), 
		(x"B631B000", x"67871DE3", x"F5DC8EF9", x"A909CBCA", x"07BE9000", x"FFF25B6C", x"4ABFD176", x"96C6828C"), 
		(x"77748000", x"39938EDB", x"A0BEB58D", x"FB3EBDDC", x"9A01A000", x"118E91EE", x"D3B8F60A", x"B5E9053A"), 
		(x"03E19000", x"63B8C8A5", x"2843A8A6", x"E5D83F4E", x"51A8A000", x"81A9A687", x"6864020D", x"651DAA5B"), 
		(x"BCDD8000", x"A9B4B9B2", x"1B62418A", x"2BCA12BD", x"253DB000", x"DB82E0F9", x"E0991F26", x"7BFB28C9"), 
		(x"C8489000", x"F39FFFCC", x"939F5CA1", x"352C902F", x"EE94B000", x"4BA5D790", x"5B45EB21", x"AB0F87A8"), 
		(x"9E5EA000", x"8DC40227", x"B1448FDA", x"C6F7B8F8", x"0D52A000", x"31C1FF3D", x"A4011E05", x"14055BFB"), 
		(x"EACBB000", x"D7EF4459", x"39B992F1", x"D8113A6A", x"C6FBA000", x"A1E6C854", x"1FDDEA02", x"C4F1F49A"), 
		(x"55F7A000", x"1DE3354E", x"0A987BDD", x"16031799", x"B26EB000", x"FBCD8E2A", x"9720F729", x"DA177608"), 
		(x"2162B000", x"47C87330", x"826566F6", x"08E5950B", x"79C7B000", x"6BEAB943", x"2CFC032E", x"0AE3D969"), 
		(x"F23CC000", x"42CB39E0", x"5AFD9229", x"94E42F6F", x"022F8000", x"CE2549E4", x"317EBCE8", x"398D5EE1"), 
		(x"86A9D000", x"18E07F9E", x"D2008F02", x"8A02ADFD", x"C9868000", x"5E027E8D", x"8AA248EF", x"E979F180"), 
		(x"3995C000", x"D2EC0E89", x"E121662E", x"4410800E", x"BD139000", x"042938F3", x"025F55C4", x"F79F7312"), 
		(x"4D00D000", x"88C748F7", x"69DC7B05", x"5AF6029C", x"76BA9000", x"940E0F9A", x"B983A1C3", x"276BDC73"), 
		(x"1B16E000", x"F69CB51C", x"4B07A87E", x"A92D2A4B", x"957C8000", x"EE6A2737", x"46C754E7", x"98610020"), 
		(x"6F83F000", x"ACB7F362", x"C3FAB555", x"B7CBA8D9", x"5ED58000", x"7E4D105E", x"FD1BA0E0", x"4895AF41"), 
		(x"D0BFE000", x"66BB8275", x"F0DB5C79", x"79D9852A", x"2A409000", x"24665620", x"75E6BDCB", x"56732DD3"), 
		(x"A42AF000", x"3C90C40B", x"78264152", x"673F07B8", x"E1E99000", x"B4416149", x"CE3A49CC", x"868782B2"), 
		(x"656FC000", x"62845733", x"2D447A26", x"350871AE", x"7C56A000", x"5A3DABCB", x"573D6EB0", x"A5A80504"), 
		(x"11FAD000", x"38AF114D", x"A5B9670D", x"2BEEF33C", x"B7FFA000", x"CA1A9CA2", x"ECE19AB7", x"755CAA65"), 
		(x"AEC6C000", x"F2A3605A", x"96988E21", x"E5FCDECF", x"C36AB000", x"9031DADC", x"641C879C", x"6BBA28F7"), 
		(x"DA53D000", x"A8882624", x"1E65930A", x"FB1A5C5D", x"08C3B000", x"0016EDB5", x"DFC0739B", x"BB4E8796"), 
		(x"8C45E000", x"D6D3DBCF", x"3CBE4071", x"08C1748A", x"EB05A000", x"7A72C518", x"208486BF", x"04445BC5"), 
		(x"F8D0F000", x"8CF89DB1", x"B4435D5A", x"1627F618", x"20ACA000", x"EA55F271", x"9B5872B8", x"D4B0F4A4"), 
		(x"47ECE000", x"46F4ECA6", x"8762B476", x"D835DBEB", x"5439B000", x"B07EB40F", x"13A56F93", x"CA567636"), 
		(x"3379F000", x"1CDFAAD8", x"0F9FA95D", x"C6D35979", x"9F90B000", x"20598366", x"A8799B94", x"1AA2D957"), 
		(x"06708000", x"526FDA2D", x"5382C538", x"4A93E323", x"1034C000", x"9532900C", x"BC847343", x"F7BB9293"), 
		(x"72E59000", x"08449C53", x"DB7FD813", x"547561B1", x"DB9DC000", x"0515A765", x"07588744", x"274F3DF2"), 
		(x"CDD98000", x"C248ED44", x"E85E313F", x"9A674C42", x"AF08D000", x"5F3EE11B", x"8FA59A6F", x"39A9BF60"), 
		(x"B94C9000", x"9863AB3A", x"60A32C14", x"8481CED0", x"64A1D000", x"CF19D672", x"34796E68", x"E95D1001"), 
		(x"EF5AA000", x"E63856D1", x"4278FF6F", x"775AE607", x"8767C000", x"B57DFEDF", x"CB3D9B4C", x"5657CC52"), 
		(x"9BCFB000", x"BC1310AF", x"CA85E244", x"69BC6495", x"4CCEC000", x"255AC9B6", x"70E16F4B", x"86A36333"), 
		(x"24F3A000", x"761F61B8", x"F9A40B68", x"A7AE4966", x"385BD000", x"7F718FC8", x"F81C7260", x"9845E1A1"), 
		(x"5066B000", x"2C3427C6", x"71591643", x"B948CBF4", x"F3F2D000", x"EF56B8A1", x"43C08667", x"48B14EC0"), 
		(x"91238000", x"7220B4FE", x"243B2D37", x"EB7FBDE2", x"6E4DE000", x"012A7223", x"DAC7A11B", x"6B9EC976"), 
		(x"E5B69000", x"280BF280", x"ACC6301C", x"F5993F70", x"A5E4E000", x"910D454A", x"611B551C", x"BB6A6617"), 
		(x"5A8A8000", x"E2078397", x"9FE7D930", x"3B8B1283", x"D171F000", x"CB260334", x"E9E64837", x"A58CE485"), 
		(x"2E1F9000", x"B82CC5E9", x"171AC41B", x"256D9011", x"1AD8F000", x"5B01345D", x"523ABC30", x"75784BE4"), 
		(x"7809A000", x"C6773802", x"35C11760", x"D6B6B8C6", x"F91EE000", x"21651CF0", x"AD7E4914", x"CA7297B7"), 
		(x"0C9CB000", x"9C5C7E7C", x"BD3C0A4B", x"C8503A54", x"32B7E000", x"B1422B99", x"16A2BD13", x"1A8638D6"), 
		(x"B3A0A000", x"56500F6B", x"8E1DE367", x"064217A7", x"4622F000", x"EB696DE7", x"9E5FA038", x"0460BA44"), 
		(x"C735B000", x"0C7B4915", x"06E0FE4C", x"18A49535", x"8D8BF000", x"7B4E5A8E", x"2583543F", x"D4941525"), 
		(x"146BC000", x"097803C5", x"DE780A93", x"84A52F51", x"F663C000", x"DE81AA29", x"3801EBF9", x"E7FA92AD"), 
		(x"60FED000", x"535345BB", x"568517B8", x"9A43ADC3", x"3DCAC000", x"4EA69D40", x"83DD1FFE", x"370E3DCC"), 
		(x"DFC2C000", x"995F34AC", x"65A4FE94", x"54518030", x"495FD000", x"148DDB3E", x"0B2002D5", x"29E8BF5E"), 
		(x"AB57D000", x"C37472D2", x"ED59E3BF", x"4AB702A2", x"82F6D000", x"84AAEC57", x"B0FCF6D2", x"F91C103F"), 
		(x"FD41E000", x"BD2F8F39", x"CF8230C4", x"B96C2A75", x"6130C000", x"FECEC4FA", x"4FB803F6", x"4616CC6C"), 
		(x"89D4F000", x"E704C947", x"477F2DEF", x"A78AA8E7", x"AA99C000", x"6EE9F393", x"F464F7F1", x"96E2630D"), 
		(x"36E8E000", x"2D08B850", x"745EC4C3", x"69988514", x"DE0CD000", x"34C2B5ED", x"7C99EADA", x"8804E19F"), 
		(x"427DF000", x"7723FE2E", x"FCA3D9E8", x"777E0786", x"15A5D000", x"A4E58284", x"C7451EDD", x"58F04EFE"), 
		(x"8338C000", x"29376D16", x"A9C1E29C", x"25497190", x"881AE000", x"4A994806", x"5E4239A1", x"7BDFC948"), 
		(x"F7ADD000", x"731C2B68", x"213CFFB7", x"3BAFF302", x"43B3E000", x"DABE7F6F", x"E59ECDA6", x"AB2B6629"), 
		(x"4891C000", x"B9105A7F", x"121D169B", x"F5BDDEF1", x"3726F000", x"80953911", x"6D63D08D", x"B5CDE4BB"), 
		(x"3C04D000", x"E33B1C01", x"9AE00BB0", x"EB5B5C63", x"FC8FF000", x"10B20E78", x"D6BF248A", x"65394BDA"), 
		(x"6A12E000", x"9D60E1EA", x"B83BD8CB", x"188074B4", x"1F49E000", x"6AD626D5", x"29FBD1AE", x"DA339789"), 
		(x"1E87F000", x"C74BA794", x"30C6C5E0", x"0666F626", x"D4E0E000", x"FAF111BC", x"922725A9", x"0AC738E8"), 
		(x"A1BBE000", x"0D47D683", x"03E72CCC", x"C874DBD5", x"A075F000", x"A0DA57C2", x"1ADA3882", x"1421BA7A"), 
		(x"D52EF000", x"576C90FD", x"8B1A31E7", x"D6925947", x"6BDCF000", x"30FD60AB", x"A106CC85", x"C4D5151B")), 
	(
		(x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000"), 
		(x"B7A40100", x"8A1F31D8", x"8589D8AB", x"E6C46464", x"734C0000", x"956FA7D6", x"A29D1297", x"6EE56854"), 
		(x"734C0000", x"956FA7D6", x"A29D1297", x"6EE56854", x"C4E80100", x"1F70960E", x"2714CA3C", x"88210C30"), 
		(x"C4E80100", x"1F70960E", x"2714CA3C", x"88210C30", x"B7A40100", x"8A1F31D8", x"8589D8AB", x"E6C46464"), 
		(x"A7B80200", x"1F128433", x"60E5F9F2", x"9E147576", x"EE260000", x"124B683E", x"80C2D68F", x"3BF3AB2C"), 
		(x"101C0300", x"950DB5EB", x"E56C2159", x"78D01112", x"9D6A0000", x"8724CFE8", x"225FC418", x"5516C378"), 
		(x"D4F40200", x"8A7D23E5", x"C278EB65", x"F0F11D22", x"2ACE0100", x"0D3BFE30", x"A7D61CB3", x"B3D2A71C"), 
		(x"63500300", x"0062123D", x"47F133CE", x"16357946", x"59820100", x"985459E6", x"054B0E24", x"DD37CF48"), 
		(x"EE260000", x"124B683E", x"80C2D68F", x"3BF3AB2C", x"499E0200", x"0D59EC0D", x"E0272F7D", x"A5E7DE5A"), 
		(x"59820100", x"985459E6", x"054B0E24", x"DD37CF48", x"3AD20200", x"98364BDB", x"42BA3DEA", x"CB02B60E"), 
		(x"9D6A0000", x"8724CFE8", x"225FC418", x"5516C378", x"8D760300", x"12297A03", x"C733E541", x"2DC6D26A"), 
		(x"2ACE0100", x"0D3BFE30", x"A7D61CB3", x"B3D2A71C", x"FE3A0300", x"8746DDD5", x"65AEF7D6", x"4323BA3E"), 
		(x"499E0200", x"0D59EC0D", x"E0272F7D", x"A5E7DE5A", x"A7B80200", x"1F128433", x"60E5F9F2", x"9E147576"), 
		(x"FE3A0300", x"8746DDD5", x"65AEF7D6", x"4323BA3E", x"D4F40200", x"8A7D23E5", x"C278EB65", x"F0F11D22"), 
		(x"3AD20200", x"98364BDB", x"42BA3DEA", x"CB02B60E", x"63500300", x"0062123D", x"47F133CE", x"16357946"), 
		(x"8D760300", x"12297A03", x"C733E541", x"2DC6D26A", x"101C0300", x"950DB5EB", x"E56C2159", x"78D01112"), 
		(x"8F3E0400", x"0D9DC877", x"6FC548E1", x"898D2CD6", x"14BD0000", x"2FBA37FF", x"6A72E5BB", x"247FEBE6"), 
		(x"389A0500", x"8782F9AF", x"EA4C904A", x"6F4948B2", x"67F10000", x"BAD59029", x"C8EFF72C", x"4A9A83B2"), 
		(x"FC720400", x"98F26FA1", x"CD585A76", x"E7684482", x"D0550100", x"30CAA1F1", x"4D662F87", x"AC5EE7D6"), 
		(x"4BD60500", x"12ED5E79", x"48D182DD", x"01AC20E6", x"A3190100", x"A5A50627", x"EFFB3D10", x"C2BB8F82"), 
		(x"28860600", x"128F4C44", x"0F20B113", x"179959A0", x"FA9B0000", x"3DF15FC1", x"EAB03334", x"1F8C40CA"), 
		(x"9F220700", x"98907D9C", x"8AA969B8", x"F15D3DC4", x"89D70000", x"A89EF817", x"482D21A3", x"7169289E"), 
		(x"5BCA0600", x"87E0EB92", x"ADBDA384", x"797C31F4", x"3E730100", x"2281C9CF", x"CDA4F908", x"97AD4CFA"), 
		(x"EC6E0700", x"0DFFDA4A", x"28347B2F", x"9FB85590", x"4D3F0100", x"B7EE6E19", x"6F39EB9F", x"F94824AE"), 
		(x"61180400", x"1FD6A049", x"EF079E6E", x"B27E87FA", x"5D230200", x"22E3DBF2", x"8A55CAC6", x"819835BC"), 
		(x"D6BC0500", x"95C99191", x"6A8E46C5", x"54BAE39E", x"2E6F0200", x"B78C7C24", x"28C8D851", x"EF7D5DE8"), 
		(x"12540400", x"8AB9079F", x"4D9A8CF9", x"DC9BEFAE", x"99CB0300", x"3D934DFC", x"AD4100FA", x"09B9398C"), 
		(x"A5F00500", x"00A63647", x"C8135452", x"3A5F8BCA", x"EA870300", x"A8FCEA2A", x"0FDC126D", x"675C51D8"), 
		(x"C6A00600", x"00C4247A", x"8FE2679C", x"2C6AF28C", x"B3050200", x"30A8B3CC", x"0A971C49", x"BA6B9E90"), 
		(x"71040700", x"8ADB15A2", x"0A6BBF37", x"CAAE96E8", x"C0490200", x"A5C7141A", x"A80A0EDE", x"D48EF6C4"), 
		(x"B5EC0600", x"95AB83AC", x"2D7F750B", x"428F9AD8", x"77ED0300", x"2FD825C2", x"2D83D675", x"324A92A0"), 
		(x"02480700", x"1FB4B274", x"A8F6ADA0", x"A44BFEBC", x"04A10300", x"BAB78214", x"8F1EC4E2", x"5CAFFAF4"), 
		(x"14BD0000", x"2FBA37FF", x"6A72E5BB", x"247FEBE6", x"9B830400", x"2227FF88", x"05B7AD5A", x"ADF2C730"), 
		(x"A3190100", x"A5A50627", x"EFFB3D10", x"C2BB8F82", x"E8CF0400", x"B748585E", x"A72ABFCD", x"C317AF64"), 
		(x"67F10000", x"BAD59029", x"C8EFF72C", x"4A9A83B2", x"5F6B0500", x"3D576986", x"22A36766", x"25D3CB00"), 
		(x"D0550100", x"30CAA1F1", x"4D662F87", x"AC5EE7D6", x"2C270500", x"A838CE50", x"803E75F1", x"4B36A354"), 
		(x"B3050200", x"30A8B3CC", x"0A971C49", x"BA6B9E90", x"75A50400", x"306C97B6", x"85757BD5", x"96016C1C"), 
		(x"04A10300", x"BAB78214", x"8F1EC4E2", x"5CAFFAF4", x"06E90400", x"A5033060", x"27E86942", x"F8E40448"), 
		(x"C0490200", x"A5C7141A", x"A80A0EDE", x"D48EF6C4", x"B14D0500", x"2F1C01B8", x"A261B1E9", x"1E20602C"), 
		(x"77ED0300", x"2FD825C2", x"2D83D675", x"324A92A0", x"C2010500", x"BA73A66E", x"00FCA37E", x"70C50878"), 
		(x"FA9B0000", x"3DF15FC1", x"EAB03334", x"1F8C40CA", x"D21D0600", x"2F7E1385", x"E5908227", x"0815196A"), 
		(x"4D3F0100", x"B7EE6E19", x"6F39EB9F", x"F94824AE", x"A1510600", x"BA11B453", x"470D90B0", x"66F0713E"), 
		(x"89D70000", x"A89EF817", x"482D21A3", x"7169289E", x"16F50700", x"300E858B", x"C284481B", x"8034155A"), 
		(x"3E730100", x"2281C9CF", x"CDA4F908", x"97AD4CFA", x"65B90700", x"A561225D", x"60195A8C", x"EED17D0E"), 
		(x"5D230200", x"22E3DBF2", x"8A55CAC6", x"819835BC", x"3C3B0600", x"3D357BBB", x"655254A8", x"33E6B246"), 
		(x"EA870300", x"A8FCEA2A", x"0FDC126D", x"675C51D8", x"4F770600", x"A85ADC6D", x"C7CF463F", x"5D03DA12"), 
		(x"2E6F0200", x"B78C7C24", x"28C8D851", x"EF7D5DE8", x"F8D30700", x"2245EDB5", x"42469E94", x"BBC7BE76"), 
		(x"99CB0300", x"3D934DFC", x"AD4100FA", x"09B9398C", x"8B9F0700", x"B72A4A63", x"E0DB8C03", x"D522D622"), 
		(x"9B830400", x"2227FF88", x"05B7AD5A", x"ADF2C730", x"8F3E0400", x"0D9DC877", x"6FC548E1", x"898D2CD6"), 
		(x"2C270500", x"A838CE50", x"803E75F1", x"4B36A354", x"FC720400", x"98F26FA1", x"CD585A76", x"E7684482"), 
		(x"E8CF0400", x"B748585E", x"A72ABFCD", x"C317AF64", x"4BD60500", x"12ED5E79", x"48D182DD", x"01AC20E6"), 
		(x"5F6B0500", x"3D576986", x"22A36766", x"25D3CB00", x"389A0500", x"8782F9AF", x"EA4C904A", x"6F4948B2"), 
		(x"3C3B0600", x"3D357BBB", x"655254A8", x"33E6B246", x"61180400", x"1FD6A049", x"EF079E6E", x"B27E87FA"), 
		(x"8B9F0700", x"B72A4A63", x"E0DB8C03", x"D522D622", x"12540400", x"8AB9079F", x"4D9A8CF9", x"DC9BEFAE"), 
		(x"4F770600", x"A85ADC6D", x"C7CF463F", x"5D03DA12", x"A5F00500", x"00A63647", x"C8135452", x"3A5F8BCA"), 
		(x"F8D30700", x"2245EDB5", x"42469E94", x"BBC7BE76", x"D6BC0500", x"95C99191", x"6A8E46C5", x"54BAE39E"), 
		(x"75A50400", x"306C97B6", x"85757BD5", x"96016C1C", x"C6A00600", x"00C4247A", x"8FE2679C", x"2C6AF28C"), 
		(x"C2010500", x"BA73A66E", x"00FCA37E", x"70C50878", x"B5EC0600", x"95AB83AC", x"2D7F750B", x"428F9AD8"), 
		(x"06E90400", x"A5033060", x"27E86942", x"F8E40448", x"02480700", x"1FB4B274", x"A8F6ADA0", x"A44BFEBC"), 
		(x"B14D0500", x"2F1C01B8", x"A261B1E9", x"1E20602C", x"71040700", x"8ADB15A2", x"0A6BBF37", x"CAAE96E8"), 
		(x"D21D0600", x"2F7E1385", x"E5908227", x"0815196A", x"28860600", x"128F4C44", x"0F20B113", x"179959A0"), 
		(x"65B90700", x"A561225D", x"60195A8C", x"EED17D0E", x"5BCA0600", x"87E0EB92", x"ADBDA384", x"797C31F4"), 
		(x"A1510600", x"BA11B453", x"470D90B0", x"66F0713E", x"EC6E0700", x"0DFFDA4A", x"28347B2F", x"9FB85590"), 
		(x"16F50700", x"300E858B", x"C284481B", x"8034155A", x"9F220700", x"98907D9C", x"8AA969B8", x"F15D3DC4"), 
		(x"DE320800", x"288350FE", x"71852AC7", x"A6BF9F96", x"E18B0000", x"5459887D", x"BF1283D3", x"1B666A73"), 
		(x"69960900", x"A29C6126", x"F40CF26C", x"407BFBF2", x"92C70000", x"C1362FAB", x"1D8F9144", x"75830227"), 
		(x"AD7E0800", x"BDECF728", x"D3183850", x"C85AF7C2", x"25630100", x"4B291E73", x"980649EF", x"93476643"), 
		(x"1ADA0900", x"37F3C6F0", x"5691E0FB", x"2E9E93A6", x"562F0100", x"DE46B9A5", x"3A9B5B78", x"FDA20E17"), 
		(x"798A0A00", x"3791D4CD", x"1160D335", x"38ABEAE0", x"0FAD0000", x"4612E043", x"3FD0555C", x"2095C15F"), 
		(x"CE2E0B00", x"BD8EE515", x"94E90B9E", x"DE6F8E84", x"7CE10000", x"D37D4795", x"9D4D47CB", x"4E70A90B"), 
		(x"0AC60A00", x"A2FE731B", x"B3FDC1A2", x"564E82B4", x"CB450100", x"5962764D", x"18C49F60", x"A8B4CD6F"), 
		(x"BD620B00", x"28E142C3", x"36741909", x"B08AE6D0", x"B8090100", x"CC0DD19B", x"BA598DF7", x"C651A53B"), 
		(x"30140800", x"3AC838C0", x"F147FC48", x"9D4C34BA", x"A8150200", x"59006470", x"5F35ACAE", x"BE81B429"), 
		(x"87B00900", x"B0D70918", x"74CE24E3", x"7B8850DE", x"DB590200", x"CC6FC3A6", x"FDA8BE39", x"D064DC7D"), 
		(x"43580800", x"AFA79F16", x"53DAEEDF", x"F3A95CEE", x"6CFD0300", x"4670F27E", x"78216692", x"36A0B819"), 
		(x"F4FC0900", x"25B8AECE", x"D6533674", x"156D388A", x"1FB10300", x"D31F55A8", x"DABC7405", x"5845D04D"), 
		(x"97AC0A00", x"25DABCF3", x"91A205BA", x"035841CC", x"46330200", x"4B4B0C4E", x"DFF77A21", x"85721F05"), 
		(x"20080B00", x"AFC58D2B", x"142BDD11", x"E59C25A8", x"357F0200", x"DE24AB98", x"7D6A68B6", x"EB977751"), 
		(x"E4E00A00", x"B0B51B25", x"333F172D", x"6DBD2998", x"82DB0300", x"543B9A40", x"F8E3B01D", x"0D531335"), 
		(x"53440B00", x"3AAA2AFD", x"B6B6CF86", x"8B794DFC", x"F1970300", x"C1543D96", x"5A7EA28A", x"63B67B61"), 
		(x"510C0C00", x"251E9889", x"1E406226", x"2F32B340", x"F5360000", x"7BE3BF82", x"D5606668", x"3F198195"), 
		(x"E6A80D00", x"AF01A951", x"9BC9BA8D", x"C9F6D724", x"867A0000", x"EE8C1854", x"77FD74FF", x"51FCE9C1"), 
		(x"22400C00", x"B0713F5F", x"BCDD70B1", x"41D7DB14", x"31DE0100", x"6493298C", x"F274AC54", x"B7388DA5"), 
		(x"95E40D00", x"3A6E0E87", x"3954A81A", x"A713BF70", x"42920100", x"F1FC8E5A", x"50E9BEC3", x"D9DDE5F1"), 
		(x"F6B40E00", x"3A0C1CBA", x"7EA59BD4", x"B126C636", x"1B100000", x"69A8D7BC", x"55A2B0E7", x"04EA2AB9"), 
		(x"41100F00", x"B0132D62", x"FB2C437F", x"57E2A252", x"685C0000", x"FCC7706A", x"F73FA270", x"6A0F42ED"), 
		(x"85F80E00", x"AF63BB6C", x"DC388943", x"DFC3AE62", x"DFF80100", x"76D841B2", x"72B67ADB", x"8CCB2689"), 
		(x"325C0F00", x"257C8AB4", x"59B151E8", x"3907CA06", x"ACB40100", x"E3B7E664", x"D02B684C", x"E22E4EDD"), 
		(x"BF2A0C00", x"3755F0B7", x"9E82B4A9", x"14C1186C", x"BCA80200", x"76BA538F", x"35474915", x"9AFE5FCF"), 
		(x"088E0D00", x"BD4AC16F", x"1B0B6C02", x"F2057C08", x"CFE40200", x"E3D5F459", x"97DA5B82", x"F41B379B"), 
		(x"CC660C00", x"A23A5761", x"3C1FA63E", x"7A247038", x"78400300", x"69CAC581", x"12538329", x"12DF53FF"), 
		(x"7BC20D00", x"282566B9", x"B9967E95", x"9CE0145C", x"0B0C0300", x"FCA56257", x"B0CE91BE", x"7C3A3BAB"), 
		(x"18920E00", x"28477484", x"FE674D5B", x"8AD56D1A", x"528E0200", x"64F13BB1", x"B5859F9A", x"A10DF4E3"), 
		(x"AF360F00", x"A258455C", x"7BEE95F0", x"6C11097E", x"21C20200", x"F19E9C67", x"17188D0D", x"CFE89CB7"), 
		(x"6BDE0E00", x"BD28D352", x"5CFA5FCC", x"E430054E", x"96660300", x"7B81ADBF", x"929155A6", x"292CF8D3"), 
		(x"DC7A0F00", x"3737E28A", x"D9738767", x"02F4612A", x"E52A0300", x"EEEE0A69", x"300C4731", x"47C99087"), 
		(x"CA8F0800", x"07396701", x"1BF7CF7C", x"82C07470", x"7A080400", x"767E77F5", x"BAA52E89", x"B694AD43"), 
		(x"7D2B0900", x"8D2656D9", x"9E7E17D7", x"64041014", x"09440400", x"E311D023", x"18383C1E", x"D871C517"), 
		(x"B9C30800", x"9256C0D7", x"B96ADDEB", x"EC251C24", x"BEE00500", x"690EE1FB", x"9DB1E4B5", x"3EB5A173"), 
		(x"0E670900", x"1849F10F", x"3CE30540", x"0AE17840", x"CDAC0500", x"FC61462D", x"3F2CF622", x"5050C927"), 
		(x"6D370A00", x"182BE332", x"7B12368E", x"1CD40106", x"942E0400", x"64351FCB", x"3A67F806", x"8D67066F"), 
		(x"DA930B00", x"9234D2EA", x"FE9BEE25", x"FA106562", x"E7620400", x"F15AB81D", x"98FAEA91", x"E3826E3B"), 
		(x"1E7B0A00", x"8D4444E4", x"D98F2419", x"72316952", x"50C60500", x"7B4589C5", x"1D73323A", x"05460A5F"), 
		(x"A9DF0B00", x"075B753C", x"5C06FCB2", x"94F50D36", x"238A0500", x"EE2A2E13", x"BFEE20AD", x"6BA3620B"), 
		(x"24A90800", x"15720F3F", x"9B3519F3", x"B933DF5C", x"33960600", x"7B279BF8", x"5A8201F4", x"13737319"), 
		(x"930D0900", x"9F6D3EE7", x"1EBCC158", x"5FF7BB38", x"40DA0600", x"EE483C2E", x"F81F1363", x"7D961B4D"), 
		(x"57E50800", x"801DA8E9", x"39A80B64", x"D7D6B708", x"F77E0700", x"64570DF6", x"7D96CBC8", x"9B527F29"), 
		(x"E0410900", x"0A029931", x"BC21D3CF", x"3112D36C", x"84320700", x"F138AA20", x"DF0BD95F", x"F5B7177D"), 
		(x"83110A00", x"0A608B0C", x"FBD0E001", x"2727AA2A", x"DDB00600", x"696CF3C6", x"DA40D77B", x"2880D835"), 
		(x"34B50B00", x"807FBAD4", x"7E5938AA", x"C1E3CE4E", x"AEFC0600", x"FC035410", x"78DDC5EC", x"4665B061"), 
		(x"F05D0A00", x"9F0F2CDA", x"594DF296", x"49C2C27E", x"19580700", x"761C65C8", x"FD541D47", x"A0A1D405"), 
		(x"47F90B00", x"15101D02", x"DCC42A3D", x"AF06A61A", x"6A140700", x"E373C21E", x"5FC90FD0", x"CE44BC51"), 
		(x"45B10C00", x"0AA4AF76", x"7432879D", x"0B4D58A6", x"6EB50400", x"59C4400A", x"D0D7CB32", x"92EB46A5"), 
		(x"F2150D00", x"80BB9EAE", x"F1BB5F36", x"ED893CC2", x"1DF90400", x"CCABE7DC", x"724AD9A5", x"FC0E2EF1"), 
		(x"36FD0C00", x"9FCB08A0", x"D6AF950A", x"65A830F2", x"AA5D0500", x"46B4D604", x"F7C3010E", x"1ACA4A95"), 
		(x"81590D00", x"15D43978", x"53264DA1", x"836C5496", x"D9110500", x"D3DB71D2", x"555E1399", x"742F22C1"), 
		(x"E2090E00", x"15B62B45", x"14D77E6F", x"95592DD0", x"80930400", x"4B8F2834", x"50151DBD", x"A918ED89"), 
		(x"55AD0F00", x"9FA91A9D", x"915EA6C4", x"739D49B4", x"F3DF0400", x"DEE08FE2", x"F2880F2A", x"C7FD85DD"), 
		(x"91450E00", x"80D98C93", x"B64A6CF8", x"FBBC4584", x"447B0500", x"54FFBE3A", x"7701D781", x"2139E1B9"), 
		(x"26E10F00", x"0AC6BD4B", x"33C3B453", x"1D7821E0", x"37370500", x"C19019EC", x"D59CC516", x"4FDC89ED"), 
		(x"AB970C00", x"18EFC748", x"F4F05112", x"30BEF38A", x"272B0600", x"549DAC07", x"30F0E44F", x"370C98FF"), 
		(x"1C330D00", x"92F0F690", x"717989B9", x"D67A97EE", x"54670600", x"C1F20BD1", x"926DF6D8", x"59E9F0AB"), 
		(x"D8DB0C00", x"8D80609E", x"566D4385", x"5E5B9BDE", x"E3C30700", x"4BED3A09", x"17E42E73", x"BF2D94CF"), 
		(x"6F7F0D00", x"079F5146", x"D3E49B2E", x"B89FFFBA", x"908F0700", x"DE829DDF", x"B5793CE4", x"D1C8FC9B"), 
		(x"0C2F0E00", x"07FD437B", x"9415A8E0", x"AEAA86FC", x"C90D0600", x"46D6C439", x"B03232C0", x"0CFF33D3"), 
		(x"BB8B0F00", x"8DE272A3", x"119C704B", x"486EE298", x"BA410600", x"D3B963EF", x"12AF2057", x"621A5B87"), 
		(x"7F630E00", x"9292E4AD", x"3688BA77", x"C04FEEA8", x"0DE50700", x"59A65237", x"9726F8FC", x"84DE3FE3"), 
		(x"C8C70F00", x"188DD575", x"B30162DC", x"268B8ACC", x"7EA90700", x"CCC9F5E1", x"35BBEA6B", x"EA3B57B7"), 
		(x"E18B0000", x"5459887D", x"BF1283D3", x"1B666A73", x"3FB90800", x"7CDAD883", x"CE97A914", x"BDD9F5E5"), 
		(x"562F0100", x"DE46B9A5", x"3A9B5B78", x"FDA20E17", x"4CF50800", x"E9B57F55", x"6C0ABB83", x"D33C9DB1"), 
		(x"92C70000", x"C1362FAB", x"1D8F9144", x"75830227", x"FB510900", x"63AA4E8D", x"E9836328", x"35F8F9D5"), 
		(x"25630100", x"4B291E73", x"980649EF", x"93476643", x"881D0900", x"F6C5E95B", x"4B1E71BF", x"5B1D9181"), 
		(x"46330200", x"4B4B0C4E", x"DFF77A21", x"85721F05", x"D19F0800", x"6E91B0BD", x"4E557F9B", x"862A5EC9"), 
		(x"F1970300", x"C1543D96", x"5A7EA28A", x"63B67B61", x"A2D30800", x"FBFE176B", x"ECC86D0C", x"E8CF369D"), 
		(x"357F0200", x"DE24AB98", x"7D6A68B6", x"EB977751", x"15770900", x"71E126B3", x"6941B5A7", x"0E0B52F9"), 
		(x"82DB0300", x"543B9A40", x"F8E3B01D", x"0D531335", x"663B0900", x"E48E8165", x"CBDCA730", x"60EE3AAD"), 
		(x"0FAD0000", x"4612E043", x"3FD0555C", x"2095C15F", x"76270A00", x"7183348E", x"2EB08669", x"183E2BBF"), 
		(x"B8090100", x"CC0DD19B", x"BA598DF7", x"C651A53B", x"056B0A00", x"E4EC9358", x"8C2D94FE", x"76DB43EB"), 
		(x"7CE10000", x"D37D4795", x"9D4D47CB", x"4E70A90B", x"B2CF0B00", x"6EF3A280", x"09A44C55", x"901F278F"), 
		(x"CB450100", x"5962764D", x"18C49F60", x"A8B4CD6F", x"C1830B00", x"FB9C0556", x"AB395EC2", x"FEFA4FDB"), 
		(x"A8150200", x"59006470", x"5F35ACAE", x"BE81B429", x"98010A00", x"63C85CB0", x"AE7250E6", x"23CD8093"), 
		(x"1FB10300", x"D31F55A8", x"DABC7405", x"5845D04D", x"EB4D0A00", x"F6A7FB66", x"0CEF4271", x"4D28E8C7"), 
		(x"DB590200", x"CC6FC3A6", x"FDA8BE39", x"D064DC7D", x"5CE90B00", x"7CB8CABE", x"89669ADA", x"ABEC8CA3"), 
		(x"6CFD0300", x"4670F27E", x"78216692", x"36A0B819", x"2FA50B00", x"E9D76D68", x"2BFB884D", x"C509E4F7"), 
		(x"6EB50400", x"59C4400A", x"D0D7CB32", x"92EB46A5", x"2B040800", x"5360EF7C", x"A4E54CAF", x"99A61E03"), 
		(x"D9110500", x"D3DB71D2", x"555E1399", x"742F22C1", x"58480800", x"C60F48AA", x"06785E38", x"F7437657"), 
		(x"1DF90400", x"CCABE7DC", x"724AD9A5", x"FC0E2EF1", x"EFEC0900", x"4C107972", x"83F18693", x"11871233"), 
		(x"AA5D0500", x"46B4D604", x"F7C3010E", x"1ACA4A95", x"9CA00900", x"D97FDEA4", x"216C9404", x"7F627A67"), 
		(x"C90D0600", x"46D6C439", x"B03232C0", x"0CFF33D3", x"C5220800", x"412B8742", x"24279A20", x"A255B52F"), 
		(x"7EA90700", x"CCC9F5E1", x"35BBEA6B", x"EA3B57B7", x"B66E0800", x"D4442094", x"86BA88B7", x"CCB0DD7B"), 
		(x"BA410600", x"D3B963EF", x"12AF2057", x"621A5B87", x"01CA0900", x"5E5B114C", x"0333501C", x"2A74B91F"), 
		(x"0DE50700", x"59A65237", x"9726F8FC", x"84DE3FE3", x"72860900", x"CB34B69A", x"A1AE428B", x"4491D14B"), 
		(x"80930400", x"4B8F2834", x"50151DBD", x"A918ED89", x"629A0A00", x"5E390371", x"44C263D2", x"3C41C059"), 
		(x"37370500", x"C19019EC", x"D59CC516", x"4FDC89ED", x"11D60A00", x"CB56A4A7", x"E65F7145", x"52A4A80D"), 
		(x"F3DF0400", x"DEE08FE2", x"F2880F2A", x"C7FD85DD", x"A6720B00", x"4149957F", x"63D6A9EE", x"B460CC69"), 
		(x"447B0500", x"54FFBE3A", x"7701D781", x"2139E1B9", x"D53E0B00", x"D42632A9", x"C14BBB79", x"DA85A43D"), 
		(x"272B0600", x"549DAC07", x"30F0E44F", x"370C98FF", x"8CBC0A00", x"4C726B4F", x"C400B55D", x"07B26B75"), 
		(x"908F0700", x"DE829DDF", x"B5793CE4", x"D1C8FC9B", x"FFF00A00", x"D91DCC99", x"669DA7CA", x"69570321"), 
		(x"54670600", x"C1F20BD1", x"926DF6D8", x"59E9F0AB", x"48540B00", x"5302FD41", x"E3147F61", x"8F936745"), 
		(x"E3C30700", x"4BED3A09", x"17E42E73", x"BF2D94CF", x"3B180B00", x"C66D5A97", x"41896DF6", x"E1760F11"), 
		(x"F5360000", x"7BE3BF82", x"D5606668", x"3F198195", x"A43A0C00", x"5EFD270B", x"CB20044E", x"102B32D5"), 
		(x"42920100", x"F1FC8E5A", x"50E9BEC3", x"D9DDE5F1", x"D7760C00", x"CB9280DD", x"69BD16D9", x"7ECE5A81"), 
		(x"867A0000", x"EE8C1854", x"77FD74FF", x"51FCE9C1", x"60D20D00", x"418DB105", x"EC34CE72", x"980A3EE5"), 
		(x"31DE0100", x"6493298C", x"F274AC54", x"B7388DA5", x"139E0D00", x"D4E216D3", x"4EA9DCE5", x"F6EF56B1"), 
		(x"528E0200", x"64F13BB1", x"B5859F9A", x"A10DF4E3", x"4A1C0C00", x"4CB64F35", x"4BE2D2C1", x"2BD899F9"), 
		(x"E52A0300", x"EEEE0A69", x"300C4731", x"47C99087", x"39500C00", x"D9D9E8E3", x"E97FC056", x"453DF1AD"), 
		(x"21C20200", x"F19E9C67", x"17188D0D", x"CFE89CB7", x"8EF40D00", x"53C6D93B", x"6CF618FD", x"A3F995C9"), 
		(x"96660300", x"7B81ADBF", x"929155A6", x"292CF8D3", x"FDB80D00", x"C6A97EED", x"CE6B0A6A", x"CD1CFD9D"), 
		(x"1B100000", x"69A8D7BC", x"55A2B0E7", x"04EA2AB9", x"EDA40E00", x"53A4CB06", x"2B072B33", x"B5CCEC8F"), 
		(x"ACB40100", x"E3B7E664", x"D02B684C", x"E22E4EDD", x"9EE80E00", x"C6CB6CD0", x"899A39A4", x"DB2984DB"), 
		(x"685C0000", x"FCC7706A", x"F73FA270", x"6A0F42ED", x"294C0F00", x"4CD45D08", x"0C13E10F", x"3DEDE0BF"), 
		(x"DFF80100", x"76D841B2", x"72B67ADB", x"8CCB2689", x"5A000F00", x"D9BBFADE", x"AE8EF398", x"530888EB"), 
		(x"BCA80200", x"76BA538F", x"35474915", x"9AFE5FCF", x"03820E00", x"41EFA338", x"ABC5FDBC", x"8E3F47A3"), 
		(x"0B0C0300", x"FCA56257", x"B0CE91BE", x"7C3A3BAB", x"70CE0E00", x"D48004EE", x"0958EF2B", x"E0DA2FF7"), 
		(x"CFE40200", x"E3D5F459", x"97DA5B82", x"F41B379B", x"C76A0F00", x"5E9F3536", x"8CD13780", x"061E4B93"), 
		(x"78400300", x"69CAC581", x"12538329", x"12DF53FF", x"B4260F00", x"CBF092E0", x"2E4C2517", x"68FB23C7"), 
		(x"7A080400", x"767E77F5", x"BAA52E89", x"B694AD43", x"B0870C00", x"714710F4", x"A152E1F5", x"3454D933"), 
		(x"CDAC0500", x"FC61462D", x"3F2CF622", x"5050C927", x"C3CB0C00", x"E428B722", x"03CFF362", x"5AB1B167"), 
		(x"09440400", x"E311D023", x"18383C1E", x"D871C517", x"746F0D00", x"6E3786FA", x"86462BC9", x"BC75D503"), 
		(x"BEE00500", x"690EE1FB", x"9DB1E4B5", x"3EB5A173", x"07230D00", x"FB58212C", x"24DB395E", x"D290BD57"), 
		(x"DDB00600", x"696CF3C6", x"DA40D77B", x"2880D835", x"5EA10C00", x"630C78CA", x"2190377A", x"0FA7721F"), 
		(x"6A140700", x"E373C21E", x"5FC90FD0", x"CE44BC51", x"2DED0C00", x"F663DF1C", x"830D25ED", x"61421A4B"), 
		(x"AEFC0600", x"FC035410", x"78DDC5EC", x"4665B061", x"9A490D00", x"7C7CEEC4", x"0684FD46", x"87867E2F"), 
		(x"19580700", x"761C65C8", x"FD541D47", x"A0A1D405", x"E9050D00", x"E9134912", x"A419EFD1", x"E963167B"), 
		(x"942E0400", x"64351FCB", x"3A67F806", x"8D67066F", x"F9190E00", x"7C1EFCF9", x"4175CE88", x"91B30769"), 
		(x"238A0500", x"EE2A2E13", x"BFEE20AD", x"6BA3620B", x"8A550E00", x"E9715B2F", x"E3E8DC1F", x"FF566F3D"), 
		(x"E7620400", x"F15AB81D", x"98FAEA91", x"E3826E3B", x"3DF10F00", x"636E6AF7", x"666104B4", x"19920B59"), 
		(x"50C60500", x"7B4589C5", x"1D73323A", x"05460A5F", x"4EBD0F00", x"F601CD21", x"C4FC1623", x"7777630D"), 
		(x"33960600", x"7B279BF8", x"5A8201F4", x"13737319", x"173F0E00", x"6E5594C7", x"C1B71807", x"AA40AC45"), 
		(x"84320700", x"F138AA20", x"DF0BD95F", x"F5B7177D", x"64730E00", x"FB3A3311", x"632A0A90", x"C4A5C411"), 
		(x"40DA0600", x"EE483C2E", x"F81F1363", x"7D961B4D", x"D3D70F00", x"712502C9", x"E6A3D23B", x"2261A075"), 
		(x"F77E0700", x"64570DF6", x"7D96CBC8", x"9B527F29", x"A09B0F00", x"E44AA51F", x"443EC0AC", x"4C84C821"), 
		(x"3FB90800", x"7CDAD883", x"CE97A914", x"BDD9F5E5", x"DE320800", x"288350FE", x"71852AC7", x"A6BF9F96"), 
		(x"881D0900", x"F6C5E95B", x"4B1E71BF", x"5B1D9181", x"AD7E0800", x"BDECF728", x"D3183850", x"C85AF7C2"), 
		(x"4CF50800", x"E9B57F55", x"6C0ABB83", x"D33C9DB1", x"1ADA0900", x"37F3C6F0", x"5691E0FB", x"2E9E93A6"), 
		(x"FB510900", x"63AA4E8D", x"E9836328", x"35F8F9D5", x"69960900", x"A29C6126", x"F40CF26C", x"407BFBF2"), 
		(x"98010A00", x"63C85CB0", x"AE7250E6", x"23CD8093", x"30140800", x"3AC838C0", x"F147FC48", x"9D4C34BA"), 
		(x"2FA50B00", x"E9D76D68", x"2BFB884D", x"C509E4F7", x"43580800", x"AFA79F16", x"53DAEEDF", x"F3A95CEE"), 
		(x"EB4D0A00", x"F6A7FB66", x"0CEF4271", x"4D28E8C7", x"F4FC0900", x"25B8AECE", x"D6533674", x"156D388A"), 
		(x"5CE90B00", x"7CB8CABE", x"89669ADA", x"ABEC8CA3", x"87B00900", x"B0D70918", x"74CE24E3", x"7B8850DE"), 
		(x"D19F0800", x"6E91B0BD", x"4E557F9B", x"862A5EC9", x"97AC0A00", x"25DABCF3", x"91A205BA", x"035841CC"), 
		(x"663B0900", x"E48E8165", x"CBDCA730", x"60EE3AAD", x"E4E00A00", x"B0B51B25", x"333F172D", x"6DBD2998"), 
		(x"A2D30800", x"FBFE176B", x"ECC86D0C", x"E8CF369D", x"53440B00", x"3AAA2AFD", x"B6B6CF86", x"8B794DFC"), 
		(x"15770900", x"71E126B3", x"6941B5A7", x"0E0B52F9", x"20080B00", x"AFC58D2B", x"142BDD11", x"E59C25A8"), 
		(x"76270A00", x"7183348E", x"2EB08669", x"183E2BBF", x"798A0A00", x"3791D4CD", x"1160D335", x"38ABEAE0"), 
		(x"C1830B00", x"FB9C0556", x"AB395EC2", x"FEFA4FDB", x"0AC60A00", x"A2FE731B", x"B3FDC1A2", x"564E82B4"), 
		(x"056B0A00", x"E4EC9358", x"8C2D94FE", x"76DB43EB", x"BD620B00", x"28E142C3", x"36741909", x"B08AE6D0"), 
		(x"B2CF0B00", x"6EF3A280", x"09A44C55", x"901F278F", x"CE2E0B00", x"BD8EE515", x"94E90B9E", x"DE6F8E84"), 
		(x"B0870C00", x"714710F4", x"A152E1F5", x"3454D933", x"CA8F0800", x"07396701", x"1BF7CF7C", x"82C07470"), 
		(x"07230D00", x"FB58212C", x"24DB395E", x"D290BD57", x"B9C30800", x"9256C0D7", x"B96ADDEB", x"EC251C24"), 
		(x"C3CB0C00", x"E428B722", x"03CFF362", x"5AB1B167", x"0E670900", x"1849F10F", x"3CE30540", x"0AE17840"), 
		(x"746F0D00", x"6E3786FA", x"86462BC9", x"BC75D503", x"7D2B0900", x"8D2656D9", x"9E7E17D7", x"64041014"), 
		(x"173F0E00", x"6E5594C7", x"C1B71807", x"AA40AC45", x"24A90800", x"15720F3F", x"9B3519F3", x"B933DF5C"), 
		(x"A09B0F00", x"E44AA51F", x"443EC0AC", x"4C84C821", x"57E50800", x"801DA8E9", x"39A80B64", x"D7D6B708"), 
		(x"64730E00", x"FB3A3311", x"632A0A90", x"C4A5C411", x"E0410900", x"0A029931", x"BC21D3CF", x"3112D36C"), 
		(x"D3D70F00", x"712502C9", x"E6A3D23B", x"2261A075", x"930D0900", x"9F6D3EE7", x"1EBCC158", x"5FF7BB38"), 
		(x"5EA10C00", x"630C78CA", x"2190377A", x"0FA7721F", x"83110A00", x"0A608B0C", x"FBD0E001", x"2727AA2A"), 
		(x"E9050D00", x"E9134912", x"A419EFD1", x"E963167B", x"F05D0A00", x"9F0F2CDA", x"594DF296", x"49C2C27E"), 
		(x"2DED0C00", x"F663DF1C", x"830D25ED", x"61421A4B", x"47F90B00", x"15101D02", x"DCC42A3D", x"AF06A61A"), 
		(x"9A490D00", x"7C7CEEC4", x"0684FD46", x"87867E2F", x"34B50B00", x"807FBAD4", x"7E5938AA", x"C1E3CE4E"), 
		(x"F9190E00", x"7C1EFCF9", x"4175CE88", x"91B30769", x"6D370A00", x"182BE332", x"7B12368E", x"1CD40106"), 
		(x"4EBD0F00", x"F601CD21", x"C4FC1623", x"7777630D", x"1E7B0A00", x"8D4444E4", x"D98F2419", x"72316952"), 
		(x"8A550E00", x"E9715B2F", x"E3E8DC1F", x"FF566F3D", x"A9DF0B00", x"075B753C", x"5C06FCB2", x"94F50D36"), 
		(x"3DF10F00", x"636E6AF7", x"666104B4", x"19920B59", x"DA930B00", x"9234D2EA", x"FE9BEE25", x"FA106562"), 
		(x"2B040800", x"5360EF7C", x"A4E54CAF", x"99A61E03", x"45B10C00", x"0AA4AF76", x"7432879D", x"0B4D58A6"), 
		(x"9CA00900", x"D97FDEA4", x"216C9404", x"7F627A67", x"36FD0C00", x"9FCB08A0", x"D6AF950A", x"65A830F2"), 
		(x"58480800", x"C60F48AA", x"06785E38", x"F7437657", x"81590D00", x"15D43978", x"53264DA1", x"836C5496"), 
		(x"EFEC0900", x"4C107972", x"83F18693", x"11871233", x"F2150D00", x"80BB9EAE", x"F1BB5F36", x"ED893CC2"), 
		(x"8CBC0A00", x"4C726B4F", x"C400B55D", x"07B26B75", x"AB970C00", x"18EFC748", x"F4F05112", x"30BEF38A"), 
		(x"3B180B00", x"C66D5A97", x"41896DF6", x"E1760F11", x"D8DB0C00", x"8D80609E", x"566D4385", x"5E5B9BDE"), 
		(x"FFF00A00", x"D91DCC99", x"669DA7CA", x"69570321", x"6F7F0D00", x"079F5146", x"D3E49B2E", x"B89FFFBA"), 
		(x"48540B00", x"5302FD41", x"E3147F61", x"8F936745", x"1C330D00", x"92F0F690", x"717989B9", x"D67A97EE"), 
		(x"C5220800", x"412B8742", x"24279A20", x"A255B52F", x"0C2F0E00", x"07FD437B", x"9415A8E0", x"AEAA86FC"), 
		(x"72860900", x"CB34B69A", x"A1AE428B", x"4491D14B", x"7F630E00", x"9292E4AD", x"3688BA77", x"C04FEEA8"), 
		(x"B66E0800", x"D4442094", x"86BA88B7", x"CCB0DD7B", x"C8C70F00", x"188DD575", x"B30162DC", x"268B8ACC"), 
		(x"01CA0900", x"5E5B114C", x"0333501C", x"2A74B91F", x"BB8B0F00", x"8DE272A3", x"119C704B", x"486EE298"), 
		(x"629A0A00", x"5E390371", x"44C263D2", x"3C41C059", x"E2090E00", x"15B62B45", x"14D77E6F", x"95592DD0"), 
		(x"D53E0B00", x"D42632A9", x"C14BBB79", x"DA85A43D", x"91450E00", x"80D98C93", x"B64A6CF8", x"FBBC4584"), 
		(x"11D60A00", x"CB56A4A7", x"E65F7145", x"52A4A80D", x"26E10F00", x"0AC6BD4B", x"33C3B453", x"1D7821E0"), 
		(x"A6720B00", x"4149957F", x"63D6A9EE", x"B460CC69", x"55AD0F00", x"9FA91A9D", x"915EA6C4", x"739D49B4"), 
		(x"A43A0C00", x"5EFD270B", x"CB20044E", x"102B32D5", x"510C0C00", x"251E9889", x"1E406226", x"2F32B340"), 
		(x"139E0D00", x"D4E216D3", x"4EA9DCE5", x"F6EF56B1", x"22400C00", x"B0713F5F", x"BCDD70B1", x"41D7DB14"), 
		(x"D7760C00", x"CB9280DD", x"69BD16D9", x"7ECE5A81", x"95E40D00", x"3A6E0E87", x"3954A81A", x"A713BF70"), 
		(x"60D20D00", x"418DB105", x"EC34CE72", x"980A3EE5", x"E6A80D00", x"AF01A951", x"9BC9BA8D", x"C9F6D724"), 
		(x"03820E00", x"41EFA338", x"ABC5FDBC", x"8E3F47A3", x"BF2A0C00", x"3755F0B7", x"9E82B4A9", x"14C1186C"), 
		(x"B4260F00", x"CBF092E0", x"2E4C2517", x"68FB23C7", x"CC660C00", x"A23A5761", x"3C1FA63E", x"7A247038"), 
		(x"70CE0E00", x"D48004EE", x"0958EF2B", x"E0DA2FF7", x"7BC20D00", x"282566B9", x"B9967E95", x"9CE0145C"), 
		(x"C76A0F00", x"5E9F3536", x"8CD13780", x"061E4B93", x"088E0D00", x"BD4AC16F", x"1B0B6C02", x"F2057C08"), 
		(x"4A1C0C00", x"4CB64F35", x"4BE2D2C1", x"2BD899F9", x"18920E00", x"28477484", x"FE674D5B", x"8AD56D1A"), 
		(x"FDB80D00", x"C6A97EED", x"CE6B0A6A", x"CD1CFD9D", x"6BDE0E00", x"BD28D352", x"5CFA5FCC", x"E430054E"), 
		(x"39500C00", x"D9D9E8E3", x"E97FC056", x"453DF1AD", x"DC7A0F00", x"3737E28A", x"D9738767", x"02F4612A"), 
		(x"8EF40D00", x"53C6D93B", x"6CF618FD", x"A3F995C9", x"AF360F00", x"A258455C", x"7BEE95F0", x"6C11097E"), 
		(x"EDA40E00", x"53A4CB06", x"2B072B33", x"B5CCEC8F", x"F6B40E00", x"3A0C1CBA", x"7EA59BD4", x"B126C636"), 
		(x"5A000F00", x"D9BBFADE", x"AE8EF398", x"530888EB", x"85F80E00", x"AF63BB6C", x"DC388943", x"DFC3AE62"), 
		(x"9EE80E00", x"C6CB6CD0", x"899A39A4", x"DB2984DB", x"325C0F00", x"257C8AB4", x"59B151E8", x"3907CA06"), 
		(x"294C0F00", x"4CD45D08", x"0C13E10F", x"3DEDE0BF", x"41100F00", x"B0132D62", x"FB2C437F", x"57E2A252")), 
	(
		(x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000"), 
		(x"515C0010", x"40F372FB", x"FCE72602", x"71575061", x"2E390000", x"64DD6689", x"3CD406FC", x"B1F490BC"), 
		(x"2E390000", x"64DD6689", x"3CD406FC", x"B1F490BC", x"7F650010", x"242E1472", x"C03320FE", x"C0A3C0DD"), 
		(x"7F650010", x"242E1472", x"C03320FE", x"C0A3C0DD", x"515C0010", x"40F372FB", x"FCE72602", x"71575061"), 
		(x"A2B80020", x"81E7E5F6", x"F9CE4C04", x"E2AFA0C0", x"5C720000", x"C9BACD12", x"79A90DF9", x"63E92178"), 
		(x"F3E40030", x"C114970D", x"05296A06", x"93F8F0A1", x"724B0000", x"AD67AB9B", x"457D0B05", x"D21DB1C4"), 
		(x"8C810020", x"E53A837F", x"C51A4AF8", x"535B307C", x"23170010", x"ED94D960", x"B99A2D07", x"A34AE1A5"), 
		(x"DDDD0030", x"A5C9F184", x"39FD6CFA", x"220C601D", x"0D2E0010", x"8949BFE9", x"854E2BFB", x"12BE7119"), 
		(x"5C720000", x"C9BACD12", x"79A90DF9", x"63E92178", x"FECA0020", x"485D28E4", x"806741FD", x"814681B8"), 
		(x"0D2E0010", x"8949BFE9", x"854E2BFB", x"12BE7119", x"D0F30020", x"2C804E6D", x"BCB34701", x"30B21104"), 
		(x"724B0000", x"AD67AB9B", x"457D0B05", x"D21DB1C4", x"81AF0030", x"6C733C96", x"40546103", x"41E54165"), 
		(x"23170010", x"ED94D960", x"B99A2D07", x"A34AE1A5", x"AF960030", x"08AE5A1F", x"7C8067FF", x"F011D1D9"), 
		(x"FECA0020", x"485D28E4", x"806741FD", x"814681B8", x"A2B80020", x"81E7E5F6", x"F9CE4C04", x"E2AFA0C0"), 
		(x"AF960030", x"08AE5A1F", x"7C8067FF", x"F011D1D9", x"8C810020", x"E53A837F", x"C51A4AF8", x"535B307C"), 
		(x"D0F30020", x"2C804E6D", x"BCB34701", x"30B21104", x"DDDD0030", x"A5C9F184", x"39FD6CFA", x"220C601D"), 
		(x"81AF0030", x"6C733C96", x"40546103", x"41E54165", x"F3E40030", x"C114970D", x"05296A06", x"93F8F0A1"), 
		(x"4DCE0040", x"3B5BEC7E", x"36656BA8", x"23633A05", x"78AB0000", x"A0CD5A34", x"5D5CA0F7", x"727784CB"), 
		(x"1C920050", x"7BA89E85", x"CA824DAA", x"52346A64", x"56920000", x"C4103CBD", x"6188A60B", x"C3831477"), 
		(x"63F70040", x"5F868AF7", x"0AB16D54", x"9297AAB9", x"07CE0010", x"84E34E46", x"9D6F8009", x"B2D44416"), 
		(x"32AB0050", x"1F75F80C", x"F6564B56", x"E3C0FAD8", x"29F70010", x"E03E28CF", x"A1BB86F5", x"0320D4AA"), 
		(x"EF760060", x"BABC0988", x"CFAB27AC", x"C1CC9AC5", x"24D90000", x"69779726", x"24F5AD0E", x"119EA5B3"), 
		(x"BE2A0070", x"FA4F7B73", x"334C01AE", x"B09BCAA4", x"0AE00000", x"0DAAF1AF", x"1821ABF2", x"A06A350F"), 
		(x"C14F0060", x"DE616F01", x"F37F2150", x"70380A79", x"5BBC0010", x"4D598354", x"E4C68DF0", x"D13D656E"), 
		(x"90130070", x"9E921DFA", x"0F980752", x"016F5A18", x"75850010", x"2984E5DD", x"D8128B0C", x"60C9F5D2"), 
		(x"11BC0040", x"F2E1216C", x"4FCC6651", x"408A1B7D", x"86610020", x"E89072D0", x"DD3BE10A", x"F3310573"), 
		(x"40E00050", x"B2125397", x"B32B4053", x"31DD4B1C", x"A8580020", x"8C4D1459", x"E1EFE7F6", x"42C595CF"), 
		(x"3F850040", x"963C47E5", x"731860AD", x"F17E8BC1", x"F9040030", x"CCBE66A2", x"1D08C1F4", x"3392C5AE"), 
		(x"6ED90050", x"D6CF351E", x"8FFF46AF", x"8029DBA0", x"D73D0030", x"A863002B", x"21DCC708", x"82665512"), 
		(x"B3040060", x"7306C49A", x"B6022A55", x"A225BBBD", x"DA130020", x"212ABFC2", x"A492ECF3", x"90D8240B"), 
		(x"E2580070", x"33F5B661", x"4AE50C57", x"D372EBDC", x"F42A0020", x"45F7D94B", x"9846EA0F", x"212CB4B7"), 
		(x"9D3D0060", x"17DBA213", x"8AD62CA9", x"13D12B01", x"A5760030", x"0504ABB0", x"64A1CC0D", x"507BE4D6"), 
		(x"CC610070", x"5728D0E8", x"76310AAB", x"62867B60", x"8B4F0030", x"61D9CD39", x"5875CAF1", x"E18F746A"), 
		(x"78AB0000", x"A0CD5A34", x"5D5CA0F7", x"727784CB", x"35650040", x"9B96B64A", x"6B39CB5F", x"5114BECE"), 
		(x"29F70010", x"E03E28CF", x"A1BB86F5", x"0320D4AA", x"1B5C0040", x"FF4BD0C3", x"57EDCDA3", x"E0E02E72"), 
		(x"56920000", x"C4103CBD", x"6188A60B", x"C3831477", x"4A000050", x"BFB8A238", x"AB0AEBA1", x"91B77E13"), 
		(x"07CE0010", x"84E34E46", x"9D6F8009", x"B2D44416", x"64390050", x"DB65C4B1", x"97DEED5D", x"2043EEAF"), 
		(x"DA130020", x"212ABFC2", x"A492ECF3", x"90D8240B", x"69170040", x"522C7B58", x"1290C6A6", x"32FD9FB6"), 
		(x"8B4F0030", x"61D9CD39", x"5875CAF1", x"E18F746A", x"472E0040", x"36F11DD1", x"2E44C05A", x"83090F0A"), 
		(x"F42A0020", x"45F7D94B", x"9846EA0F", x"212CB4B7", x"16720050", x"76026F2A", x"D2A3E658", x"F25E5F6B"), 
		(x"A5760030", x"0504ABB0", x"64A1CC0D", x"507BE4D6", x"384B0050", x"12DF09A3", x"EE77E0A4", x"43AACFD7"), 
		(x"24D90000", x"69779726", x"24F5AD0E", x"119EA5B3", x"CBAF0060", x"D3CB9EAE", x"EB5E8AA2", x"D0523F76"), 
		(x"75850010", x"2984E5DD", x"D8128B0C", x"60C9F5D2", x"E5960060", x"B716F827", x"D78A8C5E", x"61A6AFCA"), 
		(x"0AE00000", x"0DAAF1AF", x"1821ABF2", x"A06A350F", x"B4CA0070", x"F7E58ADC", x"2B6DAA5C", x"10F1FFAB"), 
		(x"5BBC0010", x"4D598354", x"E4C68DF0", x"D13D656E", x"9AF30070", x"9338EC55", x"17B9ACA0", x"A1056F17"), 
		(x"86610020", x"E89072D0", x"DD3BE10A", x"F3310573", x"97DD0060", x"1A7153BC", x"92F7875B", x"B3BB1E0E"), 
		(x"D73D0030", x"A863002B", x"21DCC708", x"82665512", x"B9E40060", x"7EAC3535", x"AE2381A7", x"024F8EB2"), 
		(x"A8580020", x"8C4D1459", x"E1EFE7F6", x"42C595CF", x"E8B80070", x"3E5F47CE", x"52C4A7A5", x"7318DED3"), 
		(x"F9040030", x"CCBE66A2", x"1D08C1F4", x"3392C5AE", x"C6810070", x"5A822147", x"6E10A159", x"C2EC4E6F"), 
		(x"35650040", x"9B96B64A", x"6B39CB5F", x"5114BECE", x"4DCE0040", x"3B5BEC7E", x"36656BA8", x"23633A05"), 
		(x"64390050", x"DB65C4B1", x"97DEED5D", x"2043EEAF", x"63F70040", x"5F868AF7", x"0AB16D54", x"9297AAB9"), 
		(x"1B5C0040", x"FF4BD0C3", x"57EDCDA3", x"E0E02E72", x"32AB0050", x"1F75F80C", x"F6564B56", x"E3C0FAD8"), 
		(x"4A000050", x"BFB8A238", x"AB0AEBA1", x"91B77E13", x"1C920050", x"7BA89E85", x"CA824DAA", x"52346A64"), 
		(x"97DD0060", x"1A7153BC", x"92F7875B", x"B3BB1E0E", x"11BC0040", x"F2E1216C", x"4FCC6651", x"408A1B7D"), 
		(x"C6810070", x"5A822147", x"6E10A159", x"C2EC4E6F", x"3F850040", x"963C47E5", x"731860AD", x"F17E8BC1"), 
		(x"B9E40060", x"7EAC3535", x"AE2381A7", x"024F8EB2", x"6ED90050", x"D6CF351E", x"8FFF46AF", x"8029DBA0"), 
		(x"E8B80070", x"3E5F47CE", x"52C4A7A5", x"7318DED3", x"40E00050", x"B2125397", x"B32B4053", x"31DD4B1C"), 
		(x"69170040", x"522C7B58", x"1290C6A6", x"32FD9FB6", x"B3040060", x"7306C49A", x"B6022A55", x"A225BBBD"), 
		(x"384B0050", x"12DF09A3", x"EE77E0A4", x"43AACFD7", x"9D3D0060", x"17DBA213", x"8AD62CA9", x"13D12B01"), 
		(x"472E0040", x"36F11DD1", x"2E44C05A", x"83090F0A", x"CC610070", x"5728D0E8", x"76310AAB", x"62867B60"), 
		(x"16720050", x"76026F2A", x"D2A3E658", x"F25E5F6B", x"E2580070", x"33F5B661", x"4AE50C57", x"D372EBDC"), 
		(x"CBAF0060", x"D3CB9EAE", x"EB5E8AA2", x"D0523F76", x"EF760060", x"BABC0988", x"CFAB27AC", x"C1CC9AC5"), 
		(x"9AF30070", x"9338EC55", x"17B9ACA0", x"A1056F17", x"C14F0060", x"DE616F01", x"F37F2150", x"70380A79"), 
		(x"E5960060", x"B716F827", x"D78A8C5E", x"61A6AFCA", x"90130070", x"9E921DFA", x"0F980752", x"016F5A18"), 
		(x"B4CA0070", x"F7E58ADC", x"2B6DAA5C", x"10F1FFAB", x"BE2A0070", x"FA4F7B73", x"334C01AE", x"B09BCAA4"), 
		(x"5BD20080", x"450F18EC", x"C2C46C55", x"F362B233", x"39A60000", x"4AB753EB", x"D14E094B", x"B772B42B"), 
		(x"0A8E0090", x"05FC6A17", x"3E234A57", x"8235E252", x"179F0000", x"2E6A3562", x"ED9A0FB7", x"06862497"), 
		(x"75EB0080", x"21D27E65", x"FE106AA9", x"4296228F", x"46C30010", x"6E994799", x"117D29B5", x"77D174F6"), 
		(x"24B70090", x"61210C9E", x"02F74CAB", x"33C172EE", x"68FA0010", x"0A442110", x"2DA92F49", x"C625E44A"), 
		(x"F96A00A0", x"C4E8FD1A", x"3B0A2051", x"11CD12F3", x"65D40000", x"830D9EF9", x"A8E704B2", x"D49B9553"), 
		(x"A83600B0", x"841B8FE1", x"C7ED0653", x"609A4292", x"4BED0000", x"E7D0F870", x"9433024E", x"656F05EF"), 
		(x"D75300A0", x"A0359B93", x"07DE26AD", x"A039824F", x"1AB10010", x"A7238A8B", x"68D4244C", x"1438558E"), 
		(x"860F00B0", x"E0C6E968", x"FB3900AF", x"D16ED22E", x"34880010", x"C3FEEC02", x"540022B0", x"A5CCC532"), 
		(x"07A00080", x"8CB5D5FE", x"BB6D61AC", x"908B934B", x"C76C0020", x"02EA7B0F", x"512948B6", x"36343593"), 
		(x"56FC0090", x"CC46A705", x"478A47AE", x"E1DCC32A", x"E9550020", x"66371D86", x"6DFD4E4A", x"87C0A52F"), 
		(x"29990080", x"E868B377", x"87B96750", x"217F03F7", x"B8090030", x"26C46F7D", x"911A6848", x"F697F54E"), 
		(x"78C50090", x"A89BC18C", x"7B5E4152", x"50285396", x"96300030", x"421909F4", x"ADCE6EB4", x"476365F2"), 
		(x"A51800A0", x"0D523008", x"42A32DA8", x"7224338B", x"9B1E0020", x"CB50B61D", x"2880454F", x"55DD14EB"), 
		(x"F44400B0", x"4DA142F3", x"BE440BAA", x"037363EA", x"B5270020", x"AF8DD094", x"145443B3", x"E4298457"), 
		(x"8B2100A0", x"698F5681", x"7E772B54", x"C3D0A337", x"E47B0030", x"EF7EA26F", x"E8B365B1", x"957ED436"), 
		(x"DA7D00B0", x"297C247A", x"82900D56", x"B287F356", x"CA420030", x"8BA3C4E6", x"D467634D", x"248A448A"), 
		(x"161C00C0", x"7E54F492", x"F4A107FD", x"D0018836", x"410D0000", x"EA7A09DF", x"8C12A9BC", x"C50530E0"), 
		(x"474000D0", x"3EA78669", x"084621FF", x"A156D857", x"6F340000", x"8EA76F56", x"B0C6AF40", x"74F1A05C"), 
		(x"382500C0", x"1A89921B", x"C8750101", x"61F5188A", x"3E680010", x"CE541DAD", x"4C218942", x"05A6F03D"), 
		(x"697900D0", x"5A7AE0E0", x"34922703", x"10A248EB", x"10510010", x"AA897B24", x"70F58FBE", x"B4526081"), 
		(x"B4A400E0", x"FFB31164", x"0D6F4BF9", x"32AE28F6", x"1D7F0000", x"23C0C4CD", x"F5BBA445", x"A6EC1198"), 
		(x"E5F800F0", x"BF40639F", x"F1886DFB", x"43F97897", x"33460000", x"471DA244", x"C96FA2B9", x"17188124"), 
		(x"9A9D00E0", x"9B6E77ED", x"31BB4D05", x"835AB84A", x"621A0010", x"07EED0BF", x"358884BB", x"664FD145"), 
		(x"CBC100F0", x"DB9D0516", x"CD5C6B07", x"F20DE82B", x"4C230010", x"6333B636", x"095C8247", x"D7BB41F9"), 
		(x"4A6E00C0", x"B7EE3980", x"8D080A04", x"B3E8A94E", x"BFC70020", x"A227213B", x"0C75E841", x"4443B158"), 
		(x"1B3200D0", x"F71D4B7B", x"71EF2C06", x"C2BFF92F", x"91FE0020", x"C6FA47B2", x"30A1EEBD", x"F5B721E4"), 
		(x"645700C0", x"D3335F09", x"B1DC0CF8", x"021C39F2", x"C0A20030", x"86093549", x"CC46C8BF", x"84E07185"), 
		(x"350B00D0", x"93C02DF2", x"4D3B2AFA", x"734B6993", x"EE9B0030", x"E2D453C0", x"F092CE43", x"3514E139"), 
		(x"E8D600E0", x"3609DC76", x"74C64600", x"5147098E", x"E3B50020", x"6B9DEC29", x"75DCE5B8", x"27AA9020"), 
		(x"B98A00F0", x"76FAAE8D", x"88216002", x"201059EF", x"CD8C0020", x"0F408AA0", x"4908E344", x"965E009C"), 
		(x"C6EF00E0", x"52D4BAFF", x"481240FC", x"E0B39932", x"9CD00030", x"4FB3F85B", x"B5EFC546", x"E70950FD"), 
		(x"97B300F0", x"1227C804", x"B4F566FE", x"91E4C953", x"B2E90030", x"2B6E9ED2", x"893BC3BA", x"56FDC041"), 
		(x"23790080", x"E5C242D8", x"9F98CCA2", x"811536F8", x"0CC30040", x"D121E5A1", x"BA77C214", x"E6660AE5"), 
		(x"72250090", x"A5313023", x"637FEAA0", x"F0426699", x"22FA0040", x"B5FC8328", x"86A3C4E8", x"57929A59"), 
		(x"0D400080", x"811F2451", x"A34CCA5E", x"30E1A644", x"73A60050", x"F50FF1D3", x"7A44E2EA", x"26C5CA38"), 
		(x"5C1C0090", x"C1EC56AA", x"5FABEC5C", x"41B6F625", x"5D9F0050", x"91D2975A", x"4690E416", x"97315A84"), 
		(x"81C100A0", x"6425A72E", x"665680A6", x"63BA9638", x"50B10040", x"189B28B3", x"C3DECFED", x"858F2B9D"), 
		(x"D09D00B0", x"24D6D5D5", x"9AB1A6A4", x"12EDC659", x"7E880040", x"7C464E3A", x"FF0AC911", x"347BBB21"), 
		(x"AFF800A0", x"00F8C1A7", x"5A82865A", x"D24E0684", x"2FD40050", x"3CB53CC1", x"03EDEF13", x"452CEB40"), 
		(x"FEA400B0", x"400BB35C", x"A665A058", x"A31956E5", x"01ED0050", x"58685A48", x"3F39E9EF", x"F4D87BFC"), 
		(x"7F0B0080", x"2C788FCA", x"E631C15B", x"E2FC1780", x"F2090060", x"997CCD45", x"3A1083E9", x"67208B5D"), 
		(x"2E570090", x"6C8BFD31", x"1AD6E759", x"93AB47E1", x"DC300060", x"FDA1ABCC", x"06C48515", x"D6D41BE1"), 
		(x"51320080", x"48A5E943", x"DAE5C7A7", x"5308873C", x"8D6C0070", x"BD52D937", x"FA23A317", x"A7834B80"), 
		(x"006E0090", x"08569BB8", x"2602E1A5", x"225FD75D", x"A3550070", x"D98FBFBE", x"C6F7A5EB", x"1677DB3C"), 
		(x"DDB300A0", x"AD9F6A3C", x"1FFF8D5F", x"0053B740", x"AE7B0060", x"50C60057", x"43B98E10", x"04C9AA25"), 
		(x"8CEF00B0", x"ED6C18C7", x"E318AB5D", x"7104E721", x"80420060", x"341B66DE", x"7F6D88EC", x"B53D3A99"), 
		(x"F38A00A0", x"C9420CB5", x"232B8BA3", x"B1A727FC", x"D11E0070", x"74E81425", x"838AAEEE", x"C46A6AF8"), 
		(x"A2D600B0", x"89B17E4E", x"DFCCADA1", x"C0F0779D", x"FF270070", x"103572AC", x"BF5EA812", x"759EFA44"), 
		(x"6EB700C0", x"DE99AEA6", x"A9FDA70A", x"A2760CFD", x"74680040", x"71ECBF95", x"E72B62E3", x"94118E2E"), 
		(x"3FEB00D0", x"9E6ADC5D", x"551A8108", x"D3215C9C", x"5A510040", x"1531D91C", x"DBFF641F", x"25E51E92"), 
		(x"408E00C0", x"BA44C82F", x"9529A1F6", x"13829C41", x"0B0D0050", x"55C2ABE7", x"2718421D", x"54B24EF3"), 
		(x"11D200D0", x"FAB7BAD4", x"69CE87F4", x"62D5CC20", x"25340050", x"311FCD6E", x"1BCC44E1", x"E546DE4F"), 
		(x"CC0F00E0", x"5F7E4B50", x"5033EB0E", x"40D9AC3D", x"281A0040", x"B8567287", x"9E826F1A", x"F7F8AF56"), 
		(x"9D5300F0", x"1F8D39AB", x"ACD4CD0C", x"318EFC5C", x"06230040", x"DC8B140E", x"A25669E6", x"460C3FEA"), 
		(x"E23600E0", x"3BA32DD9", x"6CE7EDF2", x"F12D3C81", x"577F0050", x"9C7866F5", x"5EB14FE4", x"375B6F8B"), 
		(x"B36A00F0", x"7B505F22", x"9000CBF0", x"807A6CE0", x"79460050", x"F8A5007C", x"62654918", x"86AFFF37"), 
		(x"32C500C0", x"172363B4", x"D054AAF3", x"C19F2D85", x"8AA20060", x"39B19771", x"674C231E", x"15570F96"), 
		(x"639900D0", x"57D0114F", x"2CB38CF1", x"B0C87DE4", x"A49B0060", x"5D6CF1F8", x"5B9825E2", x"A4A39F2A"), 
		(x"1CFC00C0", x"73FE053D", x"EC80AC0F", x"706BBD39", x"F5C70070", x"1D9F8303", x"A77F03E0", x"D5F4CF4B"), 
		(x"4DA000D0", x"330D77C6", x"10678A0D", x"013CED58", x"DBFE0070", x"7942E58A", x"9BAB051C", x"64005FF7"), 
		(x"907D00E0", x"96C48642", x"299AE6F7", x"23308D45", x"D6D00060", x"F00B5A63", x"1EE52EE7", x"76BE2EEE"), 
		(x"C12100F0", x"D637F4B9", x"D57DC0F5", x"5267DD24", x"F8E90060", x"94D63CEA", x"2231281B", x"C74ABE52"), 
		(x"BE4400E0", x"F219E0CB", x"154EE00B", x"92C41DF9", x"A9B50070", x"D4254E11", x"DED60E19", x"B61DEE33"), 
		(x"EF1800F0", x"B2EA9230", x"E9A9C609", x"E3934D98", x"878C0070", x"B0F82898", x"E20208E5", x"07E97E8F"), 
		(x"39A60000", x"4AB753EB", x"D14E094B", x"B772B42B", x"62740080", x"0FB84B07", x"138A651E", x"44100618"), 
		(x"68FA0010", x"0A442110", x"2DA92F49", x"C625E44A", x"4C4D0080", x"6B652D8E", x"2F5E63E2", x"F5E496A4"), 
		(x"179F0000", x"2E6A3562", x"ED9A0FB7", x"06862497", x"1D110090", x"2B965F75", x"D3B945E0", x"84B3C6C5"), 
		(x"46C30010", x"6E994799", x"117D29B5", x"77D174F6", x"33280090", x"4F4B39FC", x"EF6D431C", x"35475679"), 
		(x"9B1E0020", x"CB50B61D", x"2880454F", x"55DD14EB", x"3E060080", x"C6028615", x"6A2368E7", x"27F92760"), 
		(x"CA420030", x"8BA3C4E6", x"D467634D", x"248A448A", x"103F0080", x"A2DFE09C", x"56F76E1B", x"960DB7DC"), 
		(x"B5270020", x"AF8DD094", x"145443B3", x"E4298457", x"41630090", x"E22C9267", x"AA104819", x"E75AE7BD"), 
		(x"E47B0030", x"EF7EA26F", x"E8B365B1", x"957ED436", x"6F5A0090", x"86F1F4EE", x"96C44EE5", x"56AE7701"), 
		(x"65D40000", x"830D9EF9", x"A8E704B2", x"D49B9553", x"9CBE00A0", x"47E563E3", x"93ED24E3", x"C55687A0"), 
		(x"34880010", x"C3FEEC02", x"540022B0", x"A5CCC532", x"B28700A0", x"2338056A", x"AF39221F", x"74A2171C"), 
		(x"4BED0000", x"E7D0F870", x"9433024E", x"656F05EF", x"E3DB00B0", x"63CB7791", x"53DE041D", x"05F5477D"), 
		(x"1AB10010", x"A7238A8B", x"68D4244C", x"1438558E", x"CDE200B0", x"07161118", x"6F0A02E1", x"B401D7C1"), 
		(x"C76C0020", x"02EA7B0F", x"512948B6", x"36343593", x"C0CC00A0", x"8E5FAEF1", x"EA44291A", x"A6BFA6D8"), 
		(x"96300030", x"421909F4", x"ADCE6EB4", x"476365F2", x"EEF500A0", x"EA82C878", x"D6902FE6", x"174B3664"), 
		(x"E9550020", x"66371D86", x"6DFD4E4A", x"87C0A52F", x"BFA900B0", x"AA71BA83", x"2A7709E4", x"661C6605"), 
		(x"B8090030", x"26C46F7D", x"911A6848", x"F697F54E", x"919000B0", x"CEACDC0A", x"16A30F18", x"D7E8F6B9"), 
		(x"74680040", x"71ECBF95", x"E72B62E3", x"94118E2E", x"1ADF0080", x"AF751133", x"4ED6C5E9", x"366782D3"), 
		(x"25340050", x"311FCD6E", x"1BCC44E1", x"E546DE4F", x"34E60080", x"CBA877BA", x"7202C315", x"8793126F"), 
		(x"5A510040", x"1531D91C", x"DBFF641F", x"25E51E92", x"65BA0090", x"8B5B0541", x"8EE5E517", x"F6C4420E"), 
		(x"0B0D0050", x"55C2ABE7", x"2718421D", x"54B24EF3", x"4B830090", x"EF8663C8", x"B231E3EB", x"4730D2B2"), 
		(x"D6D00060", x"F00B5A63", x"1EE52EE7", x"76BE2EEE", x"46AD0080", x"66CFDC21", x"377FC810", x"558EA3AB"), 
		(x"878C0070", x"B0F82898", x"E20208E5", x"07E97E8F", x"68940080", x"0212BAA8", x"0BABCEEC", x"E47A3317"), 
		(x"F8E90060", x"94D63CEA", x"2231281B", x"C74ABE52", x"39C80090", x"42E1C853", x"F74CE8EE", x"952D6376"), 
		(x"A9B50070", x"D4254E11", x"DED60E19", x"B61DEE33", x"17F10090", x"263CAEDA", x"CB98EE12", x"24D9F3CA"), 
		(x"281A0040", x"B8567287", x"9E826F1A", x"F7F8AF56", x"E41500A0", x"E72839D7", x"CEB18414", x"B721036B"), 
		(x"79460050", x"F8A5007C", x"62654918", x"86AFFF37", x"CA2C00A0", x"83F55F5E", x"F26582E8", x"06D593D7"), 
		(x"06230040", x"DC8B140E", x"A25669E6", x"460C3FEA", x"9B7000B0", x"C3062DA5", x"0E82A4EA", x"7782C3B6"), 
		(x"577F0050", x"9C7866F5", x"5EB14FE4", x"375B6F8B", x"B54900B0", x"A7DB4B2C", x"3256A216", x"C676530A"), 
		(x"8AA20060", x"39B19771", x"674C231E", x"15570F96", x"B86700A0", x"2E92F4C5", x"B71889ED", x"D4C82213"), 
		(x"DBFE0070", x"7942E58A", x"9BAB051C", x"64005FF7", x"965E00A0", x"4A4F924C", x"8BCC8F11", x"653CB2AF"), 
		(x"A49B0060", x"5D6CF1F8", x"5B9825E2", x"A4A39F2A", x"C70200B0", x"0ABCE0B7", x"772BA913", x"146BE2CE"), 
		(x"F5C70070", x"1D9F8303", x"A77F03E0", x"D5F4CF4B", x"E93B00B0", x"6E61863E", x"4BFFAFEF", x"A59F7272"), 
		(x"410D0000", x"EA7A09DF", x"8C12A9BC", x"C50530E0", x"571100C0", x"942EFD4D", x"78B3AE41", x"1504B8D6"), 
		(x"10510010", x"AA897B24", x"70F58FBE", x"B4526081", x"792800C0", x"F0F39BC4", x"4467A8BD", x"A4F0286A"), 
		(x"6F340000", x"8EA76F56", x"B0C6AF40", x"74F1A05C", x"287400D0", x"B000E93F", x"B8808EBF", x"D5A7780B"), 
		(x"3E680010", x"CE541DAD", x"4C218942", x"05A6F03D", x"064D00D0", x"D4DD8FB6", x"84548843", x"6453E8B7"), 
		(x"E3B50020", x"6B9DEC29", x"75DCE5B8", x"27AA9020", x"0B6300C0", x"5D94305F", x"011AA3B8", x"76ED99AE"), 
		(x"B2E90030", x"2B6E9ED2", x"893BC3BA", x"56FDC041", x"255A00C0", x"394956D6", x"3DCEA544", x"C7190912"), 
		(x"CD8C0020", x"0F408AA0", x"4908E344", x"965E009C", x"740600D0", x"79BA242D", x"C1298346", x"B64E5973"), 
		(x"9CD00030", x"4FB3F85B", x"B5EFC546", x"E70950FD", x"5A3F00D0", x"1D6742A4", x"FDFD85BA", x"07BAC9CF"), 
		(x"1D7F0000", x"23C0C4CD", x"F5BBA445", x"A6EC1198", x"A9DB00E0", x"DC73D5A9", x"F8D4EFBC", x"9442396E"), 
		(x"4C230010", x"6333B636", x"095C8247", x"D7BB41F9", x"87E200E0", x"B8AEB320", x"C400E940", x"25B6A9D2"), 
		(x"33460000", x"471DA244", x"C96FA2B9", x"17188124", x"D6BE00F0", x"F85DC1DB", x"38E7CF42", x"54E1F9B3"), 
		(x"621A0010", x"07EED0BF", x"358884BB", x"664FD145", x"F88700F0", x"9C80A752", x"0433C9BE", x"E515690F"), 
		(x"BFC70020", x"A227213B", x"0C75E841", x"4443B158", x"F5A900E0", x"15C918BB", x"817DE245", x"F7AB1816"), 
		(x"EE9B0030", x"E2D453C0", x"F092CE43", x"3514E139", x"DB9000E0", x"71147E32", x"BDA9E4B9", x"465F88AA"), 
		(x"91FE0020", x"C6FA47B2", x"30A1EEBD", x"F5B721E4", x"8ACC00F0", x"31E70CC9", x"414EC2BB", x"3708D8CB"), 
		(x"C0A20030", x"86093549", x"CC46C8BF", x"84E07185", x"A4F500F0", x"553A6A40", x"7D9AC447", x"86FC4877"), 
		(x"0CC30040", x"D121E5A1", x"BA77C214", x"E6660AE5", x"2FBA00C0", x"34E3A779", x"25EF0EB6", x"67733C1D"), 
		(x"5D9F0050", x"91D2975A", x"4690E416", x"97315A84", x"018300C0", x"503EC1F0", x"193B084A", x"D687ACA1"), 
		(x"22FA0040", x"B5FC8328", x"86A3C4E8", x"57929A59", x"50DF00D0", x"10CDB30B", x"E5DC2E48", x"A7D0FCC0"), 
		(x"73A60050", x"F50FF1D3", x"7A44E2EA", x"26C5CA38", x"7EE600D0", x"7410D582", x"D90828B4", x"16246C7C"), 
		(x"AE7B0060", x"50C60057", x"43B98E10", x"04C9AA25", x"73C800C0", x"FD596A6B", x"5C46034F", x"049A1D65"), 
		(x"FF270070", x"103572AC", x"BF5EA812", x"759EFA44", x"5DF100C0", x"99840CE2", x"609205B3", x"B56E8DD9"), 
		(x"80420060", x"341B66DE", x"7F6D88EC", x"B53D3A99", x"0CAD00D0", x"D9777E19", x"9C7523B1", x"C439DDB8"), 
		(x"D11E0070", x"74E81425", x"838AAEEE", x"C46A6AF8", x"229400D0", x"BDAA1890", x"A0A1254D", x"75CD4D04"), 
		(x"50B10040", x"189B28B3", x"C3DECFED", x"858F2B9D", x"D17000E0", x"7CBE8F9D", x"A5884F4B", x"E635BDA5"), 
		(x"01ED0050", x"58685A48", x"3F39E9EF", x"F4D87BFC", x"FF4900E0", x"1863E914", x"995C49B7", x"57C12D19"), 
		(x"7E880040", x"7C464E3A", x"FF0AC911", x"347BBB21", x"AE1500F0", x"58909BEF", x"65BB6FB5", x"26967D78"), 
		(x"2FD40050", x"3CB53CC1", x"03EDEF13", x"452CEB40", x"802C00F0", x"3C4DFD66", x"596F6949", x"9762EDC4"), 
		(x"F2090060", x"997CCD45", x"3A1083E9", x"67208B5D", x"8D0200E0", x"B504428F", x"DC2142B2", x"85DC9CDD"), 
		(x"A3550070", x"D98FBFBE", x"C6F7A5EB", x"1677DB3C", x"A33B00E0", x"D1D92406", x"E0F5444E", x"34280C61"), 
		(x"DC300060", x"FDA1ABCC", x"06C48515", x"D6D41BE1", x"F26700F0", x"912A56FD", x"1C12624C", x"457F5C00"), 
		(x"8D6C0070", x"BD52D937", x"FA23A317", x"A7834B80", x"DC5E00F0", x"F5F73074", x"20C664B0", x"F48BCCBC"), 
		(x"62740080", x"0FB84B07", x"138A651E", x"44100618", x"5BD20080", x"450F18EC", x"C2C46C55", x"F362B233"), 
		(x"33280090", x"4F4B39FC", x"EF6D431C", x"35475679", x"75EB0080", x"21D27E65", x"FE106AA9", x"4296228F"), 
		(x"4C4D0080", x"6B652D8E", x"2F5E63E2", x"F5E496A4", x"24B70090", x"61210C9E", x"02F74CAB", x"33C172EE"), 
		(x"1D110090", x"2B965F75", x"D3B945E0", x"84B3C6C5", x"0A8E0090", x"05FC6A17", x"3E234A57", x"8235E252"), 
		(x"C0CC00A0", x"8E5FAEF1", x"EA44291A", x"A6BFA6D8", x"07A00080", x"8CB5D5FE", x"BB6D61AC", x"908B934B"), 
		(x"919000B0", x"CEACDC0A", x"16A30F18", x"D7E8F6B9", x"29990080", x"E868B377", x"87B96750", x"217F03F7"), 
		(x"EEF500A0", x"EA82C878", x"D6902FE6", x"174B3664", x"78C50090", x"A89BC18C", x"7B5E4152", x"50285396"), 
		(x"BFA900B0", x"AA71BA83", x"2A7709E4", x"661C6605", x"56FC0090", x"CC46A705", x"478A47AE", x"E1DCC32A"), 
		(x"3E060080", x"C6028615", x"6A2368E7", x"27F92760", x"A51800A0", x"0D523008", x"42A32DA8", x"7224338B"), 
		(x"6F5A0090", x"86F1F4EE", x"96C44EE5", x"56AE7701", x"8B2100A0", x"698F5681", x"7E772B54", x"C3D0A337"), 
		(x"103F0080", x"A2DFE09C", x"56F76E1B", x"960DB7DC", x"DA7D00B0", x"297C247A", x"82900D56", x"B287F356"), 
		(x"41630090", x"E22C9267", x"AA104819", x"E75AE7BD", x"F44400B0", x"4DA142F3", x"BE440BAA", x"037363EA"), 
		(x"9CBE00A0", x"47E563E3", x"93ED24E3", x"C55687A0", x"F96A00A0", x"C4E8FD1A", x"3B0A2051", x"11CD12F3"), 
		(x"CDE200B0", x"07161118", x"6F0A02E1", x"B401D7C1", x"D75300A0", x"A0359B93", x"07DE26AD", x"A039824F"), 
		(x"B28700A0", x"2338056A", x"AF39221F", x"74A2171C", x"860F00B0", x"E0C6E968", x"FB3900AF", x"D16ED22E"), 
		(x"E3DB00B0", x"63CB7791", x"53DE041D", x"05F5477D", x"A83600B0", x"841B8FE1", x"C7ED0653", x"609A4292"), 
		(x"2FBA00C0", x"34E3A779", x"25EF0EB6", x"67733C1D", x"23790080", x"E5C242D8", x"9F98CCA2", x"811536F8"), 
		(x"7EE600D0", x"7410D582", x"D90828B4", x"16246C7C", x"0D400080", x"811F2451", x"A34CCA5E", x"30E1A644"), 
		(x"018300C0", x"503EC1F0", x"193B084A", x"D687ACA1", x"5C1C0090", x"C1EC56AA", x"5FABEC5C", x"41B6F625"), 
		(x"50DF00D0", x"10CDB30B", x"E5DC2E48", x"A7D0FCC0", x"72250090", x"A5313023", x"637FEAA0", x"F0426699"), 
		(x"8D0200E0", x"B504428F", x"DC2142B2", x"85DC9CDD", x"7F0B0080", x"2C788FCA", x"E631C15B", x"E2FC1780"), 
		(x"DC5E00F0", x"F5F73074", x"20C664B0", x"F48BCCBC", x"51320080", x"48A5E943", x"DAE5C7A7", x"5308873C"), 
		(x"A33B00E0", x"D1D92406", x"E0F5444E", x"34280C61", x"006E0090", x"08569BB8", x"2602E1A5", x"225FD75D"), 
		(x"F26700F0", x"912A56FD", x"1C12624C", x"457F5C00", x"2E570090", x"6C8BFD31", x"1AD6E759", x"93AB47E1"), 
		(x"73C800C0", x"FD596A6B", x"5C46034F", x"049A1D65", x"DDB300A0", x"AD9F6A3C", x"1FFF8D5F", x"0053B740"), 
		(x"229400D0", x"BDAA1890", x"A0A1254D", x"75CD4D04", x"F38A00A0", x"C9420CB5", x"232B8BA3", x"B1A727FC"), 
		(x"5DF100C0", x"99840CE2", x"609205B3", x"B56E8DD9", x"A2D600B0", x"89B17E4E", x"DFCCADA1", x"C0F0779D"), 
		(x"0CAD00D0", x"D9777E19", x"9C7523B1", x"C439DDB8", x"8CEF00B0", x"ED6C18C7", x"E318AB5D", x"7104E721"), 
		(x"D17000E0", x"7CBE8F9D", x"A5884F4B", x"E635BDA5", x"81C100A0", x"6425A72E", x"665680A6", x"63BA9638"), 
		(x"802C00F0", x"3C4DFD66", x"596F6949", x"9762EDC4", x"AFF800A0", x"00F8C1A7", x"5A82865A", x"D24E0684"), 
		(x"FF4900E0", x"1863E914", x"995C49B7", x"57C12D19", x"FEA400B0", x"400BB35C", x"A665A058", x"A31956E5"), 
		(x"AE1500F0", x"58909BEF", x"65BB6FB5", x"26967D78", x"D09D00B0", x"24D6D5D5", x"9AB1A6A4", x"12EDC659"), 
		(x"1ADF0080", x"AF751133", x"4ED6C5E9", x"366782D3", x"6EB700C0", x"DE99AEA6", x"A9FDA70A", x"A2760CFD"), 
		(x"4B830090", x"EF8663C8", x"B231E3EB", x"4730D2B2", x"408E00C0", x"BA44C82F", x"9529A1F6", x"13829C41"), 
		(x"34E60080", x"CBA877BA", x"7202C315", x"8793126F", x"11D200D0", x"FAB7BAD4", x"69CE87F4", x"62D5CC20"), 
		(x"65BA0090", x"8B5B0541", x"8EE5E517", x"F6C4420E", x"3FEB00D0", x"9E6ADC5D", x"551A8108", x"D3215C9C"), 
		(x"B86700A0", x"2E92F4C5", x"B71889ED", x"D4C82213", x"32C500C0", x"172363B4", x"D054AAF3", x"C19F2D85"), 
		(x"E93B00B0", x"6E61863E", x"4BFFAFEF", x"A59F7272", x"1CFC00C0", x"73FE053D", x"EC80AC0F", x"706BBD39"), 
		(x"965E00A0", x"4A4F924C", x"8BCC8F11", x"653CB2AF", x"4DA000D0", x"330D77C6", x"10678A0D", x"013CED58"), 
		(x"C70200B0", x"0ABCE0B7", x"772BA913", x"146BE2CE", x"639900D0", x"57D0114F", x"2CB38CF1", x"B0C87DE4"), 
		(x"46AD0080", x"66CFDC21", x"377FC810", x"558EA3AB", x"907D00E0", x"96C48642", x"299AE6F7", x"23308D45"), 
		(x"17F10090", x"263CAEDA", x"CB98EE12", x"24D9F3CA", x"BE4400E0", x"F219E0CB", x"154EE00B", x"92C41DF9"), 
		(x"68940080", x"0212BAA8", x"0BABCEEC", x"E47A3317", x"EF1800F0", x"B2EA9230", x"E9A9C609", x"E3934D98"), 
		(x"39C80090", x"42E1C853", x"F74CE8EE", x"952D6376", x"C12100F0", x"D637F4B9", x"D57DC0F5", x"5267DD24"), 
		(x"E41500A0", x"E72839D7", x"CEB18414", x"B721036B", x"CC0F00E0", x"5F7E4B50", x"5033EB0E", x"40D9AC3D"), 
		(x"B54900B0", x"A7DB4B2C", x"3256A216", x"C676530A", x"E23600E0", x"3BA32DD9", x"6CE7EDF2", x"F12D3C81"), 
		(x"CA2C00A0", x"83F55F5E", x"F26582E8", x"06D593D7", x"B36A00F0", x"7B505F22", x"9000CBF0", x"807A6CE0"), 
		(x"9B7000B0", x"C3062DA5", x"0E82A4EA", x"7782C3B6", x"9D5300F0", x"1F8D39AB", x"ACD4CD0C", x"318EFC5C"), 
		(x"571100C0", x"942EFD4D", x"78B3AE41", x"1504B8D6", x"161C00C0", x"7E54F492", x"F4A107FD", x"D0018836"), 
		(x"064D00D0", x"D4DD8FB6", x"84548843", x"6453E8B7", x"382500C0", x"1A89921B", x"C8750101", x"61F5188A"), 
		(x"792800C0", x"F0F39BC4", x"4467A8BD", x"A4F0286A", x"697900D0", x"5A7AE0E0", x"34922703", x"10A248EB"), 
		(x"287400D0", x"B000E93F", x"B8808EBF", x"D5A7780B", x"474000D0", x"3EA78669", x"084621FF", x"A156D857"), 
		(x"F5A900E0", x"15C918BB", x"817DE245", x"F7AB1816", x"4A6E00C0", x"B7EE3980", x"8D080A04", x"B3E8A94E"), 
		(x"A4F500F0", x"553A6A40", x"7D9AC447", x"86FC4877", x"645700C0", x"D3335F09", x"B1DC0CF8", x"021C39F2"), 
		(x"DB9000E0", x"71147E32", x"BDA9E4B9", x"465F88AA", x"350B00D0", x"93C02DF2", x"4D3B2AFA", x"734B6993"), 
		(x"8ACC00F0", x"31E70CC9", x"414EC2BB", x"3708D8CB", x"1B3200D0", x"F71D4B7B", x"71EF2C06", x"C2BFF92F"), 
		(x"0B6300C0", x"5D94305F", x"011AA3B8", x"76ED99AE", x"E8D600E0", x"3609DC76", x"74C64600", x"5147098E"), 
		(x"5A3F00D0", x"1D6742A4", x"FDFD85BA", x"07BAC9CF", x"C6EF00E0", x"52D4BAFF", x"481240FC", x"E0B39932"), 
		(x"255A00C0", x"394956D6", x"3DCEA544", x"C7190912", x"97B300F0", x"1227C804", x"B4F566FE", x"91E4C953"), 
		(x"740600D0", x"79BA242D", x"C1298346", x"B64E5973", x"B98A00F0", x"76FAAE8D", x"88216002", x"201059EF"), 
		(x"A9DB00E0", x"DC73D5A9", x"F8D4EFBC", x"9442396E", x"B4A400E0", x"FFB31164", x"0D6F4BF9", x"32AE28F6"), 
		(x"F88700F0", x"9C80A752", x"0433C9BE", x"E515690F", x"9A9D00E0", x"9B6E77ED", x"31BB4D05", x"835AB84A"), 
		(x"87E200E0", x"B8AEB320", x"C400E940", x"25B6A9D2", x"CBC100F0", x"DB9D0516", x"CD5C6B07", x"F20DE82B"), 
		(x"D6BE00F0", x"F85DC1DB", x"38E7CF42", x"54E1F9B3", x"E5F800F0", x"BF40639F", x"F1886DFB", x"43F97897")), 
	(
		(x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000", x"00000000"), 
		(x"C04E0001", x"33B9C010", x"AE0EBB05", x"B5A4C63B", x"C8F10000", x"0B2DE782", x"6BF648A4", x"539CBDBF"), 
		(x"C8F10000", x"0B2DE782", x"6BF648A4", x"539CBDBF", x"08BF0001", x"38942792", x"C5F8F3A1", x"E6387B84"), 
		(x"08BF0001", x"38942792", x"C5F8F3A1", x"E6387B84", x"C04E0001", x"33B9C010", x"AE0EBB05", x"B5A4C63B"), 
		(x"88230002", x"5FE7A7B3", x"99E585AA", x"8D75F7F1", x"51AC0000", x"25E30F14", x"79E22A4C", x"1298BD46"), 
		(x"486D0003", x"6C5E67A3", x"37EB3EAF", x"38D131CA", x"995D0000", x"2ECEE896", x"121462E8", x"410400F9"), 
		(x"40D20002", x"54CA4031", x"F213CD0E", x"DEE94A4E", x"59130001", x"1D772886", x"BC1AD9ED", x"F4A0C6C2"), 
		(x"809C0003", x"67738021", x"5C1D760B", x"6B4D8C75", x"91E20001", x"165ACF04", x"D7EC9149", x"A73C7B7D"), 
		(x"51AC0000", x"25E30F14", x"79E22A4C", x"1298BD46", x"D98F0002", x"7A04A8A7", x"E007AFE6", x"9FED4AB7"), 
		(x"91E20001", x"165ACF04", x"D7EC9149", x"A73C7B7D", x"117E0002", x"71294F25", x"8BF1E742", x"CC71F708"), 
		(x"995D0000", x"2ECEE896", x"121462E8", x"410400F9", x"D1300003", x"42908F35", x"25FF5C47", x"79D53133"), 
		(x"59130001", x"1D772886", x"BC1AD9ED", x"F4A0C6C2", x"19C10003", x"49BD68B7", x"4E0914E3", x"2A498C8C"), 
		(x"D98F0002", x"7A04A8A7", x"E007AFE6", x"9FED4AB7", x"88230002", x"5FE7A7B3", x"99E585AA", x"8D75F7F1"), 
		(x"19C10003", x"49BD68B7", x"4E0914E3", x"2A498C8C", x"40D20002", x"54CA4031", x"F213CD0E", x"DEE94A4E"), 
		(x"117E0002", x"71294F25", x"8BF1E742", x"CC71F708", x"809C0003", x"67738021", x"5C1D760B", x"6B4D8C75"), 
		(x"D1300003", x"42908F35", x"25FF5C47", x"79D53133", x"486D0003", x"6C5E67A3", x"37EB3EAF", x"38D131CA"), 
		(x"D0080004", x"8C768F77", x"9DC5B050", x"AF4A29DA", x"6BA90000", x"40EBF9AA", x"98321C3D", x"76ACC733"), 
		(x"10460005", x"BFCF4F67", x"33CB0B55", x"1AEEEFE1", x"A3580000", x"4BC61E28", x"F3C45499", x"25307A8C"), 
		(x"18F90004", x"875B68F5", x"F633F8F4", x"FCD69465", x"63160001", x"787FDE38", x"5DCAEF9C", x"9094BCB7"), 
		(x"D8B70005", x"B4E2A8E5", x"583D43F1", x"4972525E", x"ABE70001", x"735239BA", x"363CA738", x"C3080108"), 
		(x"582B0006", x"D39128C4", x"042035FA", x"223FDE2B", x"3A050000", x"6508F6BE", x"E1D03671", x"64347A75"), 
		(x"98650007", x"E028E8D4", x"AA2E8EFF", x"979B1810", x"F2F40000", x"6E25113C", x"8A267ED5", x"37A8C7CA"), 
		(x"90DA0006", x"D8BCCF46", x"6FD67D5E", x"71A36394", x"32BA0001", x"5D9CD12C", x"2428C5D0", x"820C01F1"), 
		(x"50940007", x"EB050F56", x"C1D8C65B", x"C407A5AF", x"FA4B0001", x"56B136AE", x"4FDE8D74", x"D190BC4E"), 
		(x"81A40004", x"A9958063", x"E4279A1C", x"BDD2949C", x"B2260002", x"3AEF510D", x"7835B3DB", x"E9418D84"), 
		(x"41EA0005", x"9A2C4073", x"4A292119", x"087652A7", x"7AD70002", x"31C2B68F", x"13C3FB7F", x"BADD303B"), 
		(x"49550004", x"A2B867E1", x"8FD1D2B8", x"EE4E2923", x"BA990003", x"027B769F", x"BDCD407A", x"0F79F600"), 
		(x"891B0005", x"9101A7F1", x"21DF69BD", x"5BEAEF18", x"72680003", x"0956911D", x"D63B08DE", x"5CE54BBF"), 
		(x"09870006", x"F67227D0", x"7DC21FB6", x"30A7636D", x"E38A0002", x"1F0C5E19", x"01D79997", x"FBD930C2"), 
		(x"C9C90007", x"C5CBE7C0", x"D3CCA4B3", x"8503A556", x"2B7B0002", x"1421B99B", x"6A21D133", x"A8458D7D"), 
		(x"C1760006", x"FD5FC052", x"16345712", x"633BDED2", x"EB350003", x"2798798B", x"C42F6A36", x"1DE14B46"), 
		(x"01380007", x"CEE60042", x"B83AEC17", x"D69F18E9", x"23C40003", x"2CB59E09", x"AFD92292", x"4E7DF6F9"), 
		(x"6BA90000", x"40EBF9AA", x"98321C3D", x"76ACC733", x"BBA10004", x"CC9D76DD", x"05F7AC6D", x"D9E6EEE9"), 
		(x"ABE70001", x"735239BA", x"363CA738", x"C3080108", x"73500004", x"C7B0915F", x"6E01E4C9", x"8A7A5356"), 
		(x"A3580000", x"4BC61E28", x"F3C45499", x"25307A8C", x"B31E0005", x"F409514F", x"C00F5FCC", x"3FDE956D"), 
		(x"63160001", x"787FDE38", x"5DCAEF9C", x"9094BCB7", x"7BEF0005", x"FF24B6CD", x"ABF91768", x"6C4228D2"), 
		(x"E38A0002", x"1F0C5E19", x"01D79997", x"FBD930C2", x"EA0D0004", x"E97E79C9", x"7C158621", x"CB7E53AF"), 
		(x"23C40003", x"2CB59E09", x"AFD92292", x"4E7DF6F9", x"22FC0004", x"E2539E4B", x"17E3CE85", x"98E2EE10"), 
		(x"2B7B0002", x"1421B99B", x"6A21D133", x"A8458D7D", x"E2B20005", x"D1EA5E5B", x"B9ED7580", x"2D46282B"), 
		(x"EB350003", x"2798798B", x"C42F6A36", x"1DE14B46", x"2A430005", x"DAC7B9D9", x"D21B3D24", x"7EDA9594"), 
		(x"3A050000", x"6508F6BE", x"E1D03671", x"64347A75", x"622E0006", x"B699DE7A", x"E5F0038B", x"460BA45E"), 
		(x"FA4B0001", x"56B136AE", x"4FDE8D74", x"D190BC4E", x"AADF0006", x"BDB439F8", x"8E064B2F", x"159719E1"), 
		(x"F2F40000", x"6E25113C", x"8A267ED5", x"37A8C7CA", x"6A910007", x"8E0DF9E8", x"2008F02A", x"A033DFDA"), 
		(x"32BA0001", x"5D9CD12C", x"2428C5D0", x"820C01F1", x"A2600007", x"85201E6A", x"4BFEB88E", x"F3AF6265"), 
		(x"B2260002", x"3AEF510D", x"7835B3DB", x"E9418D84", x"33820006", x"937AD16E", x"9C1229C7", x"54931918"), 
		(x"72680003", x"0956911D", x"D63B08DE", x"5CE54BBF", x"FB730006", x"985736EC", x"F7E46163", x"070FA4A7"), 
		(x"7AD70002", x"31C2B68F", x"13C3FB7F", x"BADD303B", x"3B3D0007", x"ABEEF6FC", x"59EADA66", x"B2AB629C"), 
		(x"BA990003", x"027B769F", x"BDCD407A", x"0F79F600", x"F3CC0007", x"A0C3117E", x"321C92C2", x"E137DF23"), 
		(x"BBA10004", x"CC9D76DD", x"05F7AC6D", x"D9E6EEE9", x"D0080004", x"8C768F77", x"9DC5B050", x"AF4A29DA"), 
		(x"7BEF0005", x"FF24B6CD", x"ABF91768", x"6C4228D2", x"18F90004", x"875B68F5", x"F633F8F4", x"FCD69465"), 
		(x"73500004", x"C7B0915F", x"6E01E4C9", x"8A7A5356", x"D8B70005", x"B4E2A8E5", x"583D43F1", x"4972525E"), 
		(x"B31E0005", x"F409514F", x"C00F5FCC", x"3FDE956D", x"10460005", x"BFCF4F67", x"33CB0B55", x"1AEEEFE1"), 
		(x"33820006", x"937AD16E", x"9C1229C7", x"54931918", x"81A40004", x"A9958063", x"E4279A1C", x"BDD2949C"), 
		(x"F3CC0007", x"A0C3117E", x"321C92C2", x"E137DF23", x"49550004", x"A2B867E1", x"8FD1D2B8", x"EE4E2923"), 
		(x"FB730006", x"985736EC", x"F7E46163", x"070FA4A7", x"891B0005", x"9101A7F1", x"21DF69BD", x"5BEAEF18"), 
		(x"3B3D0007", x"ABEEF6FC", x"59EADA66", x"B2AB629C", x"41EA0005", x"9A2C4073", x"4A292119", x"087652A7"), 
		(x"EA0D0004", x"E97E79C9", x"7C158621", x"CB7E53AF", x"09870006", x"F67227D0", x"7DC21FB6", x"30A7636D"), 
		(x"2A430005", x"DAC7B9D9", x"D21B3D24", x"7EDA9594", x"C1760006", x"FD5FC052", x"16345712", x"633BDED2"), 
		(x"22FC0004", x"E2539E4B", x"17E3CE85", x"98E2EE10", x"01380007", x"CEE60042", x"B83AEC17", x"D69F18E9"), 
		(x"E2B20005", x"D1EA5E5B", x"B9ED7580", x"2D46282B", x"C9C90007", x"C5CBE7C0", x"D3CCA4B3", x"8503A556"), 
		(x"622E0006", x"B699DE7A", x"E5F0038B", x"460BA45E", x"582B0006", x"D39128C4", x"042035FA", x"223FDE2B"), 
		(x"A2600007", x"85201E6A", x"4BFEB88E", x"F3AF6265", x"90DA0006", x"D8BCCF46", x"6FD67D5E", x"71A36394"), 
		(x"AADF0006", x"BDB439F8", x"8E064B2F", x"159719E1", x"50940007", x"EB050F56", x"C1D8C65B", x"C407A5AF"), 
		(x"6A910007", x"8E0DF9E8", x"2008F02A", x"A033DFDA", x"98650007", x"E028E8D4", x"AA2E8EFF", x"979B1810"), 
		(x"A8AE0008", x"2079397D", x"FE739301", x"B8A92831", x"171C0000", x"B26E3344", x"9E6A837E", x"58F8485F"), 
		(x"68E00009", x"13C0F96D", x"507D2804", x"0D0DEE0A", x"DFED0000", x"B943D4C6", x"F59CCBDA", x"0B64F5E0"), 
		(x"605F0008", x"2B54DEFF", x"9585DBA5", x"EB35958E", x"1FA30001", x"8AFA14D6", x"5B9270DF", x"BEC033DB"), 
		(x"A0110009", x"18ED1EEF", x"3B8B60A0", x"5E9153B5", x"D7520001", x"81D7F354", x"3064387B", x"ED5C8E64"), 
		(x"208D000A", x"7F9E9ECE", x"679616AB", x"35DCDFC0", x"46B00000", x"978D3C50", x"E788A932", x"4A60F519"), 
		(x"E0C3000B", x"4C275EDE", x"C998ADAE", x"807819FB", x"8E410000", x"9CA0DBD2", x"8C7EE196", x"19FC48A6"), 
		(x"E87C000A", x"74B3794C", x"0C605E0F", x"6640627F", x"4E0F0001", x"AF191BC2", x"22705A93", x"AC588E9D"), 
		(x"2832000B", x"470AB95C", x"A26EE50A", x"D3E4A444", x"86FE0001", x"A434FC40", x"49861237", x"FFC43322"), 
		(x"F9020008", x"059A3669", x"8791B94D", x"AA319577", x"CE930002", x"C86A9BE3", x"7E6D2C98", x"C71502E8"), 
		(x"394C0009", x"3623F679", x"299F0248", x"1F95534C", x"06620002", x"C3477C61", x"159B643C", x"9489BF57"), 
		(x"31F30008", x"0EB7D1EB", x"EC67F1E9", x"F9AD28C8", x"C62C0003", x"F0FEBC71", x"BB95DF39", x"212D796C"), 
		(x"F1BD0009", x"3D0E11FB", x"42694AEC", x"4C09EEF3", x"0EDD0003", x"FBD35BF3", x"D063979D", x"72B1C4D3"), 
		(x"7121000A", x"5A7D91DA", x"1E743CE7", x"27446286", x"9F3F0002", x"ED8994F7", x"078F06D4", x"D58DBFAE"), 
		(x"B16F000B", x"69C451CA", x"B07A87E2", x"92E0A4BD", x"57CE0002", x"E6A47375", x"6C794E70", x"86110211"), 
		(x"B9D0000A", x"51507658", x"75827443", x"74D8DF39", x"97800003", x"D51DB365", x"C277F575", x"33B5C42A"), 
		(x"799E000B", x"62E9B648", x"DB8CCF46", x"C17C1902", x"5F710003", x"DE3054E7", x"A981BDD1", x"60297995"), 
		(x"78A6000C", x"AC0FB60A", x"63B62351", x"17E301EB", x"7CB50000", x"F285CAEE", x"06589F43", x"2E548F6C"), 
		(x"B8E8000D", x"9FB6761A", x"CDB89854", x"A247C7D0", x"B4440000", x"F9A82D6C", x"6DAED7E7", x"7DC832D3"), 
		(x"B057000C", x"A7225188", x"08406BF5", x"447FBC54", x"740A0001", x"CA11ED7C", x"C3A06CE2", x"C86CF4E8"), 
		(x"7019000D", x"949B9198", x"A64ED0F0", x"F1DB7A6F", x"BCFB0001", x"C13C0AFE", x"A8562446", x"9BF04957"), 
		(x"F085000E", x"F3E811B9", x"FA53A6FB", x"9A96F61A", x"2D190000", x"D766C5FA", x"7FBAB50F", x"3CCC322A"), 
		(x"30CB000F", x"C051D1A9", x"545D1DFE", x"2F323021", x"E5E80000", x"DC4B2278", x"144CFDAB", x"6F508F95"), 
		(x"3874000E", x"F8C5F63B", x"91A5EE5F", x"C90A4BA5", x"25A60001", x"EFF2E268", x"BA4246AE", x"DAF449AE"), 
		(x"F83A000F", x"CB7C362B", x"3FAB555A", x"7CAE8D9E", x"ED570001", x"E4DF05EA", x"D1B40E0A", x"8968F411"), 
		(x"290A000C", x"89ECB91E", x"1A54091D", x"057BBCAD", x"A53A0002", x"88816249", x"E65F30A5", x"B1B9C5DB"), 
		(x"E944000D", x"BA55790E", x"B45AB218", x"B0DF7A96", x"6DCB0002", x"83AC85CB", x"8DA97801", x"E2257864"), 
		(x"E1FB000C", x"82C15E9C", x"71A241B9", x"56E70112", x"AD850003", x"B01545DB", x"23A7C304", x"5781BE5F"), 
		(x"21B5000D", x"B1789E8C", x"DFACFABC", x"E343C729", x"65740003", x"BB38A259", x"48518BA0", x"041D03E0"), 
		(x"A129000E", x"D60B1EAD", x"83B18CB7", x"880E4B5C", x"F4960002", x"AD626D5D", x"9FBD1AE9", x"A321789D"), 
		(x"6167000F", x"E5B2DEBD", x"2DBF37B2", x"3DAA8D67", x"3C670002", x"A64F8ADF", x"F44B524D", x"F0BDC522"), 
		(x"69D8000E", x"DD26F92F", x"E847C413", x"DB92F6E3", x"FC290003", x"95F64ACF", x"5A45E948", x"45190319"), 
		(x"A996000F", x"EE9F393F", x"46497F16", x"6E3630D8", x"34D80003", x"9EDBAD4D", x"31B3A1EC", x"1685BEA6"), 
		(x"C3070008", x"6092C0D7", x"66418F3C", x"CE05EF02", x"ACBD0004", x"7EF34599", x"9B9D2F13", x"811EA6B6"), 
		(x"03490009", x"532B00C7", x"C84F3439", x"7BA12939", x"644C0004", x"75DEA21B", x"F06B67B7", x"D2821B09"), 
		(x"0BF60008", x"6BBF2755", x"0DB7C798", x"9D9952BD", x"A4020005", x"4667620B", x"5E65DCB2", x"6726DD32"), 
		(x"CBB80009", x"5806E745", x"A3B97C9D", x"283D9486", x"6CF30005", x"4D4A8589", x"35939416", x"34BA608D"), 
		(x"4B24000A", x"3F756764", x"FFA40A96", x"437018F3", x"FD110004", x"5B104A8D", x"E27F055F", x"93861BF0"), 
		(x"8B6A000B", x"0CCCA774", x"51AAB193", x"F6D4DEC8", x"35E00004", x"503DAD0F", x"89894DFB", x"C01AA64F"), 
		(x"83D5000A", x"345880E6", x"94524232", x"10ECA54C", x"F5AE0005", x"63846D1F", x"2787F6FE", x"75BE6074"), 
		(x"439B000B", x"07E140F6", x"3A5CF937", x"A5486377", x"3D5F0005", x"68A98A9D", x"4C71BE5A", x"2622DDCB"), 
		(x"92AB0008", x"4571CFC3", x"1FA3A570", x"DC9D5244", x"75320006", x"04F7ED3E", x"7B9A80F5", x"1EF3EC01"), 
		(x"52E50009", x"76C80FD3", x"B1AD1E75", x"6939947F", x"BDC30006", x"0FDA0ABC", x"106CC851", x"4D6F51BE"), 
		(x"5A5A0008", x"4E5C2841", x"7455EDD4", x"8F01EFFB", x"7D8D0007", x"3C63CAAC", x"BE627354", x"F8CB9785"), 
		(x"9A140009", x"7DE5E851", x"DA5B56D1", x"3AA529C0", x"B57C0007", x"374E2D2E", x"D5943BF0", x"AB572A3A"), 
		(x"1A88000A", x"1A966870", x"864620DA", x"51E8A5B5", x"249E0006", x"2114E22A", x"0278AAB9", x"0C6B5147"), 
		(x"DAC6000B", x"292FA860", x"28489BDF", x"E44C638E", x"EC6F0006", x"2A3905A8", x"698EE21D", x"5FF7ECF8"), 
		(x"D279000A", x"11BB8FF2", x"EDB0687E", x"0274180A", x"2C210007", x"1980C5B8", x"C7805918", x"EA532AC3"), 
		(x"1237000B", x"22024FE2", x"43BED37B", x"B7D0DE31", x"E4D00007", x"12AD223A", x"AC7611BC", x"B9CF977C"), 
		(x"130F000C", x"ECE44FA0", x"FB843F6C", x"614FC6D8", x"C7140004", x"3E18BC33", x"03AF332E", x"F7B26185"), 
		(x"D341000D", x"DF5D8FB0", x"558A8469", x"D4EB00E3", x"0FE50004", x"35355BB1", x"68597B8A", x"A42EDC3A"), 
		(x"DBFE000C", x"E7C9A822", x"907277C8", x"32D37B67", x"CFAB0005", x"068C9BA1", x"C657C08F", x"118A1A01"), 
		(x"1BB0000D", x"D4706832", x"3E7CCCCD", x"8777BD5C", x"075A0005", x"0DA17C23", x"ADA1882B", x"4216A7BE"), 
		(x"9B2C000E", x"B303E813", x"6261BAC6", x"EC3A3129", x"96B80004", x"1BFBB327", x"7A4D1962", x"E52ADCC3"), 
		(x"5B62000F", x"80BA2803", x"CC6F01C3", x"599EF712", x"5E490004", x"10D654A5", x"11BB51C6", x"B6B6617C"), 
		(x"53DD000E", x"B82E0F91", x"0997F262", x"BFA68C96", x"9E070005", x"236F94B5", x"BFB5EAC3", x"0312A747"), 
		(x"9393000F", x"8B97CF81", x"A7994967", x"0A024AAD", x"56F60005", x"28427337", x"D443A267", x"508E1AF8"), 
		(x"42A3000C", x"C90740B4", x"82661520", x"73D77B9E", x"1E9B0006", x"441C1494", x"E3A89CC8", x"685F2B32"), 
		(x"82ED000D", x"FABE80A4", x"2C68AE25", x"C673BDA5", x"D66A0006", x"4F31F316", x"885ED46C", x"3BC3968D"), 
		(x"8A52000C", x"C22AA736", x"E9905D84", x"204BC621", x"16240007", x"7C883306", x"26506F69", x"8E6750B6"), 
		(x"4A1C000D", x"F1936726", x"479EE681", x"95EF001A", x"DED50007", x"77A5D484", x"4DA627CD", x"DDFBED09"), 
		(x"CA80000E", x"96E0E707", x"1B83908A", x"FEA28C6F", x"4F370006", x"61FF1B80", x"9A4AB684", x"7AC79674"), 
		(x"0ACE000F", x"A5592717", x"B58D2B8F", x"4B064A54", x"87C60006", x"6AD2FC02", x"F1BCFE20", x"295B2BCB"), 
		(x"0271000E", x"9DCD0085", x"7075D82E", x"AD3E31D0", x"47880007", x"596B3C12", x"5FB24525", x"9CFFEDF0"), 
		(x"C23F000F", x"AE74C095", x"DE7B632B", x"189AF7EB", x"8F790007", x"5246DB90", x"34440D81", x"CF63504F"), 
		(x"171C0000", x"B26E3344", x"9E6A837E", x"58F8485F", x"BFB20008", x"92170A39", x"6019107F", x"E051606E"), 
		(x"D7520001", x"81D7F354", x"3064387B", x"ED5C8E64", x"77430008", x"993AEDBB", x"0BEF58DB", x"B3CDDDD1"), 
		(x"DFED0000", x"B943D4C6", x"F59CCBDA", x"0B64F5E0", x"B70D0009", x"AA832DAB", x"A5E1E3DE", x"06691BEA"), 
		(x"1FA30001", x"8AFA14D6", x"5B9270DF", x"BEC033DB", x"7FFC0009", x"A1AECA29", x"CE17AB7A", x"55F5A655"), 
		(x"9F3F0002", x"ED8994F7", x"078F06D4", x"D58DBFAE", x"EE1E0008", x"B7F4052D", x"19FB3A33", x"F2C9DD28"), 
		(x"5F710003", x"DE3054E7", x"A981BDD1", x"60297995", x"26EF0008", x"BCD9E2AF", x"720D7297", x"A1556097"), 
		(x"57CE0002", x"E6A47375", x"6C794E70", x"86110211", x"E6A10009", x"8F6022BF", x"DC03C992", x"14F1A6AC"), 
		(x"97800003", x"D51DB365", x"C277F575", x"33B5C42A", x"2E500009", x"844DC53D", x"B7F58136", x"476D1B13"), 
		(x"46B00000", x"978D3C50", x"E788A932", x"4A60F519", x"663D000A", x"E813A29E", x"801EBF99", x"7FBC2AD9"), 
		(x"86FE0001", x"A434FC40", x"49861237", x"FFC43322", x"AECC000A", x"E33E451C", x"EBE8F73D", x"2C209766"), 
		(x"8E410000", x"9CA0DBD2", x"8C7EE196", x"19FC48A6", x"6E82000B", x"D087850C", x"45E64C38", x"9984515D"), 
		(x"4E0F0001", x"AF191BC2", x"22705A93", x"AC588E9D", x"A673000B", x"DBAA628E", x"2E10049C", x"CA18ECE2"), 
		(x"CE930002", x"C86A9BE3", x"7E6D2C98", x"C71502E8", x"3791000A", x"CDF0AD8A", x"F9FC95D5", x"6D24979F"), 
		(x"0EDD0003", x"FBD35BF3", x"D063979D", x"72B1C4D3", x"FF60000A", x"C6DD4A08", x"920ADD71", x"3EB82A20"), 
		(x"06620002", x"C3477C61", x"159B643C", x"9489BF57", x"3F2E000B", x"F5648A18", x"3C046674", x"8B1CEC1B"), 
		(x"C62C0003", x"F0FEBC71", x"BB95DF39", x"212D796C", x"F7DF000B", x"FE496D9A", x"57F22ED0", x"D88051A4"), 
		(x"C7140004", x"3E18BC33", x"03AF332E", x"F7B26185", x"D41B0008", x"D2FCF393", x"F82B0C42", x"96FDA75D"), 
		(x"075A0005", x"0DA17C23", x"ADA1882B", x"4216A7BE", x"1CEA0008", x"D9D11411", x"93DD44E6", x"C5611AE2"), 
		(x"0FE50004", x"35355BB1", x"68597B8A", x"A42EDC3A", x"DCA40009", x"EA68D401", x"3DD3FFE3", x"70C5DCD9"), 
		(x"CFAB0005", x"068C9BA1", x"C657C08F", x"118A1A01", x"14550009", x"E1453383", x"5625B747", x"23596166"), 
		(x"4F370006", x"61FF1B80", x"9A4AB684", x"7AC79674", x"85B70008", x"F71FFC87", x"81C9260E", x"84651A1B"), 
		(x"8F790007", x"5246DB90", x"34440D81", x"CF63504F", x"4D460008", x"FC321B05", x"EA3F6EAA", x"D7F9A7A4"), 
		(x"87C60006", x"6AD2FC02", x"F1BCFE20", x"295B2BCB", x"8D080009", x"CF8BDB15", x"4431D5AF", x"625D619F"), 
		(x"47880007", x"596B3C12", x"5FB24525", x"9CFFEDF0", x"45F90009", x"C4A63C97", x"2FC79D0B", x"31C1DC20"), 
		(x"96B80004", x"1BFBB327", x"7A4D1962", x"E52ADCC3", x"0D94000A", x"A8F85B34", x"182CA3A4", x"0910EDEA"), 
		(x"56F60005", x"28427337", x"D443A267", x"508E1AF8", x"C565000A", x"A3D5BCB6", x"73DAEB00", x"5A8C5055"), 
		(x"5E490004", x"10D654A5", x"11BB51C6", x"B6B6617C", x"052B000B", x"906C7CA6", x"DDD45005", x"EF28966E"), 
		(x"9E070005", x"236F94B5", x"BFB5EAC3", x"0312A747", x"CDDA000B", x"9B419B24", x"B62218A1", x"BCB42BD1"), 
		(x"1E9B0006", x"441C1494", x"E3A89CC8", x"685F2B32", x"5C38000A", x"8D1B5420", x"61CE89E8", x"1B8850AC"), 
		(x"DED50007", x"77A5D484", x"4DA627CD", x"DDFBED09", x"94C9000A", x"8636B3A2", x"0A38C14C", x"4814ED13"), 
		(x"D66A0006", x"4F31F316", x"885ED46C", x"3BC3968D", x"5487000B", x"B58F73B2", x"A4367A49", x"FDB02B28"), 
		(x"16240007", x"7C883306", x"26506F69", x"8E6750B6", x"9C76000B", x"BEA29430", x"CFC032ED", x"AE2C9697"), 
		(x"7CB50000", x"F285CAEE", x"06589F43", x"2E548F6C", x"0413000C", x"5E8A7CE4", x"65EEBC12", x"39B78E87"), 
		(x"BCFB0001", x"C13C0AFE", x"A8562446", x"9BF04957", x"CCE2000C", x"55A79B66", x"0E18F4B6", x"6A2B3338"), 
		(x"B4440000", x"F9A82D6C", x"6DAED7E7", x"7DC832D3", x"0CAC000D", x"661E5B76", x"A0164FB3", x"DF8FF503"), 
		(x"740A0001", x"CA11ED7C", x"C3A06CE2", x"C86CF4E8", x"C45D000D", x"6D33BCF4", x"CBE00717", x"8C1348BC"), 
		(x"F4960002", x"AD626D5D", x"9FBD1AE9", x"A321789D", x"55BF000C", x"7B6973F0", x"1C0C965E", x"2B2F33C1"), 
		(x"34D80003", x"9EDBAD4D", x"31B3A1EC", x"1685BEA6", x"9D4E000C", x"70449472", x"77FADEFA", x"78B38E7E"), 
		(x"3C670002", x"A64F8ADF", x"F44B524D", x"F0BDC522", x"5D00000D", x"43FD5462", x"D9F465FF", x"CD174845"), 
		(x"FC290003", x"95F64ACF", x"5A45E948", x"45190319", x"95F1000D", x"48D0B3E0", x"B2022D5B", x"9E8BF5FA"), 
		(x"2D190000", x"D766C5FA", x"7FBAB50F", x"3CCC322A", x"DD9C000E", x"248ED443", x"85E913F4", x"A65AC430"), 
		(x"ED570001", x"E4DF05EA", x"D1B40E0A", x"8968F411", x"156D000E", x"2FA333C1", x"EE1F5B50", x"F5C6798F"), 
		(x"E5E80000", x"DC4B2278", x"144CFDAB", x"6F508F95", x"D523000F", x"1C1AF3D1", x"4011E055", x"4062BFB4"), 
		(x"25A60001", x"EFF2E268", x"BA4246AE", x"DAF449AE", x"1DD2000F", x"17371453", x"2BE7A8F1", x"13FE020B"), 
		(x"A53A0002", x"88816249", x"E65F30A5", x"B1B9C5DB", x"8C30000E", x"016DDB57", x"FC0B39B8", x"B4C27976"), 
		(x"65740003", x"BB38A259", x"48518BA0", x"041D03E0", x"44C1000E", x"0A403CD5", x"97FD711C", x"E75EC4C9"), 
		(x"6DCB0002", x"83AC85CB", x"8DA97801", x"E2257864", x"848F000F", x"39F9FCC5", x"39F3CA19", x"52FA02F2"), 
		(x"AD850003", x"B01545DB", x"23A7C304", x"5781BE5F", x"4C7E000F", x"32D41B47", x"520582BD", x"0166BF4D"), 
		(x"ACBD0004", x"7EF34599", x"9B9D2F13", x"811EA6B6", x"6FBA000C", x"1E61854E", x"FDDCA02F", x"4F1B49B4"), 
		(x"6CF30005", x"4D4A8589", x"35939416", x"34BA608D", x"A74B000C", x"154C62CC", x"962AE88B", x"1C87F40B"), 
		(x"644C0004", x"75DEA21B", x"F06B67B7", x"D2821B09", x"6705000D", x"26F5A2DC", x"3824538E", x"A9233230"), 
		(x"A4020005", x"4667620B", x"5E65DCB2", x"6726DD32", x"AFF4000D", x"2DD8455E", x"53D21B2A", x"FABF8F8F"), 
		(x"249E0006", x"2114E22A", x"0278AAB9", x"0C6B5147", x"3E16000C", x"3B828A5A", x"843E8A63", x"5D83F4F2"), 
		(x"E4D00007", x"12AD223A", x"AC7611BC", x"B9CF977C", x"F6E7000C", x"30AF6DD8", x"EFC8C2C7", x"0E1F494D"), 
		(x"EC6F0006", x"2A3905A8", x"698EE21D", x"5FF7ECF8", x"36A9000D", x"0316ADC8", x"41C679C2", x"BBBB8F76"), 
		(x"2C210007", x"1980C5B8", x"C7805918", x"EA532AC3", x"FE58000D", x"083B4A4A", x"2A303166", x"E82732C9"), 
		(x"FD110004", x"5B104A8D", x"E27F055F", x"93861BF0", x"B635000E", x"64652DE9", x"1DDB0FC9", x"D0F60303"), 
		(x"3D5F0005", x"68A98A9D", x"4C71BE5A", x"2622DDCB", x"7EC4000E", x"6F48CA6B", x"762D476D", x"836ABEBC"), 
		(x"35E00004", x"503DAD0F", x"89894DFB", x"C01AA64F", x"BE8A000F", x"5CF10A7B", x"D823FC68", x"36CE7887"), 
		(x"F5AE0005", x"63846D1F", x"2787F6FE", x"75BE6074", x"767B000F", x"57DCEDF9", x"B3D5B4CC", x"6552C538"), 
		(x"75320006", x"04F7ED3E", x"7B9A80F5", x"1EF3EC01", x"E799000E", x"418622FD", x"64392585", x"C26EBE45"), 
		(x"B57C0007", x"374E2D2E", x"D5943BF0", x"AB572A3A", x"2F68000E", x"4AABC57F", x"0FCF6D21", x"91F203FA"), 
		(x"BDC30006", x"0FDA0ABC", x"106CC851", x"4D6F51BE", x"EF26000F", x"7912056F", x"A1C1D624", x"2456C5C1"), 
		(x"7D8D0007", x"3C63CAAC", x"BE627354", x"F8CB9785", x"27D7000F", x"723FE2ED", x"CA379E80", x"77CA787E"), 
		(x"BFB20008", x"92170A39", x"6019107F", x"E051606E", x"A8AE0008", x"2079397D", x"FE739301", x"B8A92831"), 
		(x"7FFC0009", x"A1AECA29", x"CE17AB7A", x"55F5A655", x"605F0008", x"2B54DEFF", x"9585DBA5", x"EB35958E"), 
		(x"77430008", x"993AEDBB", x"0BEF58DB", x"B3CDDDD1", x"A0110009", x"18ED1EEF", x"3B8B60A0", x"5E9153B5"), 
		(x"B70D0009", x"AA832DAB", x"A5E1E3DE", x"06691BEA", x"68E00009", x"13C0F96D", x"507D2804", x"0D0DEE0A"), 
		(x"3791000A", x"CDF0AD8A", x"F9FC95D5", x"6D24979F", x"F9020008", x"059A3669", x"8791B94D", x"AA319577"), 
		(x"F7DF000B", x"FE496D9A", x"57F22ED0", x"D88051A4", x"31F30008", x"0EB7D1EB", x"EC67F1E9", x"F9AD28C8"), 
		(x"FF60000A", x"C6DD4A08", x"920ADD71", x"3EB82A20", x"F1BD0009", x"3D0E11FB", x"42694AEC", x"4C09EEF3"), 
		(x"3F2E000B", x"F5648A18", x"3C046674", x"8B1CEC1B", x"394C0009", x"3623F679", x"299F0248", x"1F95534C"), 
		(x"EE1E0008", x"B7F4052D", x"19FB3A33", x"F2C9DD28", x"7121000A", x"5A7D91DA", x"1E743CE7", x"27446286"), 
		(x"2E500009", x"844DC53D", x"B7F58136", x"476D1B13", x"B9D0000A", x"51507658", x"75827443", x"74D8DF39"), 
		(x"26EF0008", x"BCD9E2AF", x"720D7297", x"A1556097", x"799E000B", x"62E9B648", x"DB8CCF46", x"C17C1902"), 
		(x"E6A10009", x"8F6022BF", x"DC03C992", x"14F1A6AC", x"B16F000B", x"69C451CA", x"B07A87E2", x"92E0A4BD"), 
		(x"663D000A", x"E813A29E", x"801EBF99", x"7FBC2AD9", x"208D000A", x"7F9E9ECE", x"679616AB", x"35DCDFC0"), 
		(x"A673000B", x"DBAA628E", x"2E10049C", x"CA18ECE2", x"E87C000A", x"74B3794C", x"0C605E0F", x"6640627F"), 
		(x"AECC000A", x"E33E451C", x"EBE8F73D", x"2C209766", x"2832000B", x"470AB95C", x"A26EE50A", x"D3E4A444"), 
		(x"6E82000B", x"D087850C", x"45E64C38", x"9984515D", x"E0C3000B", x"4C275EDE", x"C998ADAE", x"807819FB"), 
		(x"6FBA000C", x"1E61854E", x"FDDCA02F", x"4F1B49B4", x"C3070008", x"6092C0D7", x"66418F3C", x"CE05EF02"), 
		(x"AFF4000D", x"2DD8455E", x"53D21B2A", x"FABF8F8F", x"0BF60008", x"6BBF2755", x"0DB7C798", x"9D9952BD"), 
		(x"A74B000C", x"154C62CC", x"962AE88B", x"1C87F40B", x"CBB80009", x"5806E745", x"A3B97C9D", x"283D9486"), 
		(x"6705000D", x"26F5A2DC", x"3824538E", x"A9233230", x"03490009", x"532B00C7", x"C84F3439", x"7BA12939"), 
		(x"E799000E", x"418622FD", x"64392585", x"C26EBE45", x"92AB0008", x"4571CFC3", x"1FA3A570", x"DC9D5244"), 
		(x"27D7000F", x"723FE2ED", x"CA379E80", x"77CA787E", x"5A5A0008", x"4E5C2841", x"7455EDD4", x"8F01EFFB"), 
		(x"2F68000E", x"4AABC57F", x"0FCF6D21", x"91F203FA", x"9A140009", x"7DE5E851", x"DA5B56D1", x"3AA529C0"), 
		(x"EF26000F", x"7912056F", x"A1C1D624", x"2456C5C1", x"52E50009", x"76C80FD3", x"B1AD1E75", x"6939947F"), 
		(x"3E16000C", x"3B828A5A", x"843E8A63", x"5D83F4F2", x"1A88000A", x"1A966870", x"864620DA", x"51E8A5B5"), 
		(x"FE58000D", x"083B4A4A", x"2A303166", x"E82732C9", x"D279000A", x"11BB8FF2", x"EDB0687E", x"0274180A"), 
		(x"F6E7000C", x"30AF6DD8", x"EFC8C2C7", x"0E1F494D", x"1237000B", x"22024FE2", x"43BED37B", x"B7D0DE31"), 
		(x"36A9000D", x"0316ADC8", x"41C679C2", x"BBBB8F76", x"DAC6000B", x"292FA860", x"28489BDF", x"E44C638E"), 
		(x"B635000E", x"64652DE9", x"1DDB0FC9", x"D0F60303", x"4B24000A", x"3F756764", x"FFA40A96", x"437018F3"), 
		(x"767B000F", x"57DCEDF9", x"B3D5B4CC", x"6552C538", x"83D5000A", x"345880E6", x"94524232", x"10ECA54C"), 
		(x"7EC4000E", x"6F48CA6B", x"762D476D", x"836ABEBC", x"439B000B", x"07E140F6", x"3A5CF937", x"A5486377"), 
		(x"BE8A000F", x"5CF10A7B", x"D823FC68", x"36CE7887", x"8B6A000B", x"0CCCA774", x"51AAB193", x"F6D4DEC8"), 
		(x"D41B0008", x"D2FCF393", x"F82B0C42", x"96FDA75D", x"130F000C", x"ECE44FA0", x"FB843F6C", x"614FC6D8"), 
		(x"14550009", x"E1453383", x"5625B747", x"23596166", x"DBFE000C", x"E7C9A822", x"907277C8", x"32D37B67"), 
		(x"1CEA0008", x"D9D11411", x"93DD44E6", x"C5611AE2", x"1BB0000D", x"D4706832", x"3E7CCCCD", x"8777BD5C"), 
		(x"DCA40009", x"EA68D401", x"3DD3FFE3", x"70C5DCD9", x"D341000D", x"DF5D8FB0", x"558A8469", x"D4EB00E3"), 
		(x"5C38000A", x"8D1B5420", x"61CE89E8", x"1B8850AC", x"42A3000C", x"C90740B4", x"82661520", x"73D77B9E"), 
		(x"9C76000B", x"BEA29430", x"CFC032ED", x"AE2C9697", x"8A52000C", x"C22AA736", x"E9905D84", x"204BC621"), 
		(x"94C9000A", x"8636B3A2", x"0A38C14C", x"4814ED13", x"4A1C000D", x"F1936726", x"479EE681", x"95EF001A"), 
		(x"5487000B", x"B58F73B2", x"A4367A49", x"FDB02B28", x"82ED000D", x"FABE80A4", x"2C68AE25", x"C673BDA5"), 
		(x"85B70008", x"F71FFC87", x"81C9260E", x"84651A1B", x"CA80000E", x"96E0E707", x"1B83908A", x"FEA28C6F"), 
		(x"45F90009", x"C4A63C97", x"2FC79D0B", x"31C1DC20", x"0271000E", x"9DCD0085", x"7075D82E", x"AD3E31D0"), 
		(x"4D460008", x"FC321B05", x"EA3F6EAA", x"D7F9A7A4", x"C23F000F", x"AE74C095", x"DE7B632B", x"189AF7EB"), 
		(x"8D080009", x"CF8BDB15", x"4431D5AF", x"625D619F", x"0ACE000F", x"A5592717", x"B58D2B8F", x"4B064A54"), 
		(x"0D94000A", x"A8F85B34", x"182CA3A4", x"0910EDEA", x"9B2C000E", x"B303E813", x"6261BAC6", x"EC3A3129"), 
		(x"CDDA000B", x"9B419B24", x"B62218A1", x"BCB42BD1", x"53DD000E", x"B82E0F91", x"0997F262", x"BFA68C96"), 
		(x"C565000A", x"A3D5BCB6", x"73DAEB00", x"5A8C5055", x"9393000F", x"8B97CF81", x"A7994967", x"0A024AAD"), 
		(x"052B000B", x"906C7CA6", x"DDD45005", x"EF28966E", x"5B62000F", x"80BA2803", x"CC6F01C3", x"599EF712"), 
		(x"0413000C", x"5E8A7CE4", x"65EEBC12", x"39B78E87", x"78A6000C", x"AC0FB60A", x"63B62351", x"17E301EB"), 
		(x"C45D000D", x"6D33BCF4", x"CBE00717", x"8C1348BC", x"B057000C", x"A7225188", x"08406BF5", x"447FBC54"), 
		(x"CCE2000C", x"55A79B66", x"0E18F4B6", x"6A2B3338", x"7019000D", x"949B9198", x"A64ED0F0", x"F1DB7A6F"), 
		(x"0CAC000D", x"661E5B76", x"A0164FB3", x"DF8FF503", x"B8E8000D", x"9FB6761A", x"CDB89854", x"A247C7D0"), 
		(x"8C30000E", x"016DDB57", x"FC0B39B8", x"B4C27976", x"290A000C", x"89ECB91E", x"1A54091D", x"057BBCAD"), 
		(x"4C7E000F", x"32D41B47", x"520582BD", x"0166BF4D", x"E1FB000C", x"82C15E9C", x"71A241B9", x"56E70112"), 
		(x"44C1000E", x"0A403CD5", x"97FD711C", x"E75EC4C9", x"21B5000D", x"B1789E8C", x"DFACFABC", x"E343C729"), 
		(x"848F000F", x"39F9FCC5", x"39F3CA19", x"52FA02F2", x"E944000D", x"BA55790E", x"B45AB218", x"B0DF7A96"), 
		(x"55BF000C", x"7B6973F0", x"1C0C965E", x"2B2F33C1", x"A129000E", x"D60B1EAD", x"83B18CB7", x"880E4B5C"), 
		(x"95F1000D", x"48D0B3E0", x"B2022D5B", x"9E8BF5FA", x"69D8000E", x"DD26F92F", x"E847C413", x"DB92F6E3"), 
		(x"9D4E000C", x"70449472", x"77FADEFA", x"78B38E7E", x"A996000F", x"EE9F393F", x"46497F16", x"6E3630D8"), 
		(x"5D00000D", x"43FD5462", x"D9F465FF", x"CD174845", x"6167000F", x"E5B2DEBD", x"2DBF37B2", x"3DAA8D67"), 
		(x"DD9C000E", x"248ED443", x"85E913F4", x"A65AC430", x"F085000E", x"F3E811B9", x"FA53A6FB", x"9A96F61A"), 
		(x"1DD2000F", x"17371453", x"2BE7A8F1", x"13FE020B", x"3874000E", x"F8C5F63B", x"91A5EE5F", x"C90A4BA5"), 
		(x"156D000E", x"2FA333C1", x"EE1F5B50", x"F5C6798F", x"F83A000F", x"CB7C362B", x"3FAB555A", x"7CAE8D9E"), 
		(x"D523000F", x"1C1AF3D1", x"4011E055", x"4062BFB4", x"30CB000F", x"C051D1A9", x"545D1DFE", x"2F323021"))
	);
end package;