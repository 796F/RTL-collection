library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
use ieee.std_logic_textio.all;

package blakePkg is

  constant WWIDTH : integer := 64;      -- WORD WIDTH
  constant NROUND : integer := 16;      -- ROUND NUMBER

  -----------------------------------------------------------------------------
  -- c Constants
  -----------------------------------------------------------------------------
  type c_const is array (0 to 15) of std_logic_vector(63 downto 0);  

  constant C  : c_const := ((x"243F6A8885A308D3"), (x"13198A2E03707344"),
                            (x"A4093822299F31D0"), (x"082EFA98EC4E6C89"),
                            (x"452821E638D01377"), (x"BE5466CF34E90C6C"),
                            (x"C0AC29B7C97C50DD"), (x"3F84D5B5B5470917"),
                            (x"9216D5D98979FB1B"), (x"D1310BA698DFB5AC"),
                            (x"2FFD72DBD01ADFB7"), (x"B8E1AFED6A267E96"),
                            (x"BA7C9045F12C7F99"), (x"24A19947B3916CF7"),
                            (x"0801F2E2858EFC16"), (x"636920D871574E69"));


  -----------------------------------------------------------------------------
  -- o Permutations
  -----------------------------------------------------------------------------
  type perm is array (0 to 9, 0 to 15) of integer;
  
  constant PMATRIX : perm := ((0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15),
                              (14, 10, 4, 8, 9, 15, 13, 6, 1, 12, 0, 2, 11, 7, 5, 3),
                              (11, 8, 12, 0, 5, 2, 15, 13, 10, 14, 3, 6, 7, 1, 9, 4),
                              (7, 9, 3, 1, 13, 12, 11, 14, 2, 6, 5, 10, 4, 0, 15, 8),
                              (9, 0, 5, 7, 2, 4, 10, 15, 14, 1, 11, 12, 6, 8, 3, 13),
                              (2, 12, 6, 10, 0, 11, 8, 3, 4, 13, 7, 5, 15, 14, 1, 9),
                              (12, 5, 1, 15, 14, 13, 4, 10, 0, 7, 6, 3, 9, 2, 8, 11),
                              (13, 11, 7, 14, 12, 1, 3, 9, 5, 0, 15, 4, 8, 6, 2, 10),
                              (6, 15, 14, 9, 11, 3, 0, 8, 12, 2, 13, 7, 1, 4, 10, 5),
                              (10, 2, 8, 4, 7, 6, 1, 5, 15, 11, 9, 14, 3, 12, 13, 0));

  -----------------------------------------------------------------------------
  -- i Iterations
  -----------------------------------------------------------------------------
  type iter is array (0 to 7, 0 to 3) of integer;
  
  constant IMATRIX : iter := ((0, 4, 8, 12), (1, 5, 9, 13), (2, 6, 10, 14), (3, 7, 11, 15),
                              (0, 5, 10, 15), (1, 6, 11, 12), (2, 7, 8, 13), (3, 4, 9, 14));

  
end blakePkg;
