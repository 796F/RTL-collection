//////////////////////////////////////////////////////////////////////////
//2010 CESCA @ Virginia Tech
//////////////////////////////////////////////////////////////////////////
//This program is free software: you can redistribute it and/or modify
//it under the terms of the GNU General Public License as published by
//the Free Software Foundation, either version 3 of the License, or
//(at your option) any later version.
//
//This program is distributed in the hope that it will be useful,
//but WITHOUT ANY WARRANTY; without even the implied warranty of
//MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//GNU General Public License for more details.
//
//You should have received a copy of the GNU General Public License
//along with this program.  If not, see <http://www.gnu.org/licenses/>.
//////////////////////////////////////////////////////////////////////////
module TABLE0(
	           byte_in,
	           table_out);

input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'hc04e0001
	         : (byte_in == 8'h02)? 32'hc8f10000
	         : (byte_in == 8'h03)? 32'h08bf0001
	         : (byte_in == 8'h04)? 32'h88230002
	         : (byte_in == 8'h05)? 32'h486d0003
	         : (byte_in == 8'h06)? 32'h40d20002
	         : (byte_in == 8'h07)? 32'h809c0003
	         : (byte_in == 8'h08)? 32'h51ac0000
	         : (byte_in == 8'h09)? 32'h91e20001
	         : (byte_in == 8'h0a)? 32'h995d0000
	         : (byte_in == 8'h0b)? 32'h59130001
	         : (byte_in == 8'h0c)? 32'hd98f0002
	         : (byte_in == 8'h0d)? 32'h19c10003
	         : (byte_in == 8'h0e)? 32'h117e0002
	         : (byte_in == 8'h0f)? 32'hd1300003
	         : (byte_in == 8'h10)? 32'hd0080004
	         : (byte_in == 8'h11)? 32'h10460005
	         : (byte_in == 8'h12)? 32'h18f90004
	         : (byte_in == 8'h13)? 32'hd8b70005
	         : (byte_in == 8'h14)? 32'h582b0006
	         : (byte_in == 8'h15)? 32'h98650007
	         : (byte_in == 8'h16)? 32'h90da0006
	         : (byte_in == 8'h17)? 32'h50940007
	         : (byte_in == 8'h18)? 32'h81a40004
	         : (byte_in == 8'h19)? 32'h41ea0005
	         : (byte_in == 8'h1a)? 32'h49550004
	         : (byte_in == 8'h1b)? 32'h891b0005
	         : (byte_in == 8'h1c)? 32'h09870006
	         : (byte_in == 8'h1d)? 32'hc9c90007
	         : (byte_in == 8'h1e)? 32'hc1760006
	         : (byte_in == 8'h1f)? 32'h01380007
	         : (byte_in == 8'h20)? 32'h6ba90000
	         : (byte_in == 8'h21)? 32'habe70001
	         : (byte_in == 8'h22)? 32'ha3580000
	         : (byte_in == 8'h23)? 32'h63160001
	         : (byte_in == 8'h24)? 32'he38a0002
	         : (byte_in == 8'h25)? 32'h23c40003
	         : (byte_in == 8'h26)? 32'h2b7b0002
	         : (byte_in == 8'h27)? 32'heb350003
	         : (byte_in == 8'h28)? 32'h3a050000
	         : (byte_in == 8'h29)? 32'hfa4b0001
	         : (byte_in == 8'h2a)? 32'hf2f40000
	         : (byte_in == 8'h2b)? 32'h32ba0001
	         : (byte_in == 8'h2c)? 32'hb2260002
	         : (byte_in == 8'h2d)? 32'h72680003
	         : (byte_in == 8'h2e)? 32'h7ad70002
	         : (byte_in == 8'h2f)? 32'hba990003
	         : (byte_in == 8'h30)? 32'hbba10004
	         : (byte_in == 8'h31)? 32'h7bef0005
	         : (byte_in == 8'h32)? 32'h73500004
	         : (byte_in == 8'h33)? 32'hb31e0005
	         : (byte_in == 8'h34)? 32'h33820006
	         : (byte_in == 8'h35)? 32'hf3cc0007
	         : (byte_in == 8'h36)? 32'hfb730006
	         : (byte_in == 8'h37)? 32'h3b3d0007
	         : (byte_in == 8'h38)? 32'hea0d0004
	         : (byte_in == 8'h39)? 32'h2a430005
	         : (byte_in == 8'h3a)? 32'h22fc0004
	         : (byte_in == 8'h3b)? 32'he2b20005
	         : (byte_in == 8'h3c)? 32'h622e0006
	         : (byte_in == 8'h3d)? 32'ha2600007
	         : (byte_in == 8'h3e)? 32'haadf0006
	         : (byte_in == 8'h3f)? 32'h6a910007
	         : (byte_in == 8'h40)? 32'ha8ae0008
	         : (byte_in == 8'h41)? 32'h68e00009
	         : (byte_in == 8'h42)? 32'h605f0008
	         : (byte_in == 8'h43)? 32'ha0110009
	         : (byte_in == 8'h44)? 32'h208d000a
	         : (byte_in == 8'h45)? 32'he0c3000b
	         : (byte_in == 8'h46)? 32'he87c000a
	         : (byte_in == 8'h47)? 32'h2832000b
	         : (byte_in == 8'h48)? 32'hf9020008
	         : (byte_in == 8'h49)? 32'h394c0009
	         : (byte_in == 8'h4a)? 32'h31f30008
	         : (byte_in == 8'h4b)? 32'hf1bd0009
	         : (byte_in == 8'h4c)? 32'h7121000a
	         : (byte_in == 8'h4d)? 32'hb16f000b
	         : (byte_in == 8'h4e)? 32'hb9d0000a
	         : (byte_in == 8'h4f)? 32'h799e000b
	         : (byte_in == 8'h50)? 32'h78a6000c
	         : (byte_in == 8'h51)? 32'hb8e8000d
	         : (byte_in == 8'h52)? 32'hb057000c
	         : (byte_in == 8'h53)? 32'h7019000d
	         : (byte_in == 8'h54)? 32'hf085000e
	         : (byte_in == 8'h55)? 32'h30cb000f
	         : (byte_in == 8'h56)? 32'h3874000e
	         : (byte_in == 8'h57)? 32'hf83a000f
	         : (byte_in == 8'h58)? 32'h290a000c
	         : (byte_in == 8'h59)? 32'he944000d
	         : (byte_in == 8'h5a)? 32'he1fb000c
	         : (byte_in == 8'h5b)? 32'h21b5000d
	         : (byte_in == 8'h5c)? 32'ha129000e
	         : (byte_in == 8'h5d)? 32'h6167000f
	         : (byte_in == 8'h5e)? 32'h69d8000e
	         : (byte_in == 8'h5f)? 32'ha996000f
	         : (byte_in == 8'h60)? 32'hc3070008
	         : (byte_in == 8'h61)? 32'h03490009
	         : (byte_in == 8'h62)? 32'h0bf60008
	         : (byte_in == 8'h63)? 32'hcbb80009
	         : (byte_in == 8'h64)? 32'h4b24000a
	         : (byte_in == 8'h65)? 32'h8b6a000b
	         : (byte_in == 8'h66)? 32'h83d5000a
	         : (byte_in == 8'h67)? 32'h439b000b
	         : (byte_in == 8'h68)? 32'h92ab0008
	         : (byte_in == 8'h69)? 32'h52e50009
	         : (byte_in == 8'h6a)? 32'h5a5a0008
	         : (byte_in == 8'h6b)? 32'h9a140009
	         : (byte_in == 8'h6c)? 32'h1a88000a
	         : (byte_in == 8'h6d)? 32'hdac6000b
	         : (byte_in == 8'h6e)? 32'hd279000a
	         : (byte_in == 8'h6f)? 32'h1237000b
	         : (byte_in == 8'h70)? 32'h130f000c
	         : (byte_in == 8'h71)? 32'hd341000d
	         : (byte_in == 8'h72)? 32'hdbfe000c
	         : (byte_in == 8'h73)? 32'h1bb0000d
	         : (byte_in == 8'h74)? 32'h9b2c000e
	         : (byte_in == 8'h75)? 32'h5b62000f
	         : (byte_in == 8'h76)? 32'h53dd000e
	         : (byte_in == 8'h77)? 32'h9393000f
	         : (byte_in == 8'h78)? 32'h42a3000c
	         : (byte_in == 8'h79)? 32'h82ed000d
	         : (byte_in == 8'h7a)? 32'h8a52000c
	         : (byte_in == 8'h7b)? 32'h4a1c000d
	         : (byte_in == 8'h7c)? 32'hca80000e
	         : (byte_in == 8'h7d)? 32'h0ace000f
	         : (byte_in == 8'h7e)? 32'h0271000e
	         : (byte_in == 8'h7f)? 32'hc23f000f
	         : (byte_in == 8'h80)? 32'h171c0000
	         : (byte_in == 8'h81)? 32'hd7520001
	         : (byte_in == 8'h82)? 32'hdfed0000
	         : (byte_in == 8'h83)? 32'h1fa30001
	         : (byte_in == 8'h84)? 32'h9f3f0002
	         : (byte_in == 8'h85)? 32'h5f710003
	         : (byte_in == 8'h86)? 32'h57ce0002
	         : (byte_in == 8'h87)? 32'h97800003
	         : (byte_in == 8'h88)? 32'h46b00000
	         : (byte_in == 8'h89)? 32'h86fe0001
	         : (byte_in == 8'h8a)? 32'h8e410000
	         : (byte_in == 8'h8b)? 32'h4e0f0001
	         : (byte_in == 8'h8c)? 32'hce930002
	         : (byte_in == 8'h8d)? 32'h0edd0003
	         : (byte_in == 8'h8e)? 32'h06620002
	         : (byte_in == 8'h8f)? 32'hc62c0003
	         : (byte_in == 8'h90)? 32'hc7140004
	         : (byte_in == 8'h91)? 32'h075a0005
	         : (byte_in == 8'h92)? 32'h0fe50004
	         : (byte_in == 8'h93)? 32'hcfab0005
	         : (byte_in == 8'h94)? 32'h4f370006
	         : (byte_in == 8'h95)? 32'h8f790007
	         : (byte_in == 8'h96)? 32'h87c60006
	         : (byte_in == 8'h97)? 32'h47880007
	         : (byte_in == 8'h98)? 32'h96b80004
	         : (byte_in == 8'h99)? 32'h56f60005
	         : (byte_in == 8'h9a)? 32'h5e490004
	         : (byte_in == 8'h9b)? 32'h9e070005
	         : (byte_in == 8'h9c)? 32'h1e9b0006
	         : (byte_in == 8'h9d)? 32'hded50007
	         : (byte_in == 8'h9e)? 32'hd66a0006
	         : (byte_in == 8'h9f)? 32'h16240007
	         : (byte_in == 8'ha0)? 32'h7cb50000
	         : (byte_in == 8'ha1)? 32'hbcfb0001
	         : (byte_in == 8'ha2)? 32'hb4440000
	         : (byte_in == 8'ha3)? 32'h740a0001
	         : (byte_in == 8'ha4)? 32'hf4960002
	         : (byte_in == 8'ha5)? 32'h34d80003
	         : (byte_in == 8'ha6)? 32'h3c670002
	         : (byte_in == 8'ha7)? 32'hfc290003
	         : (byte_in == 8'ha8)? 32'h2d190000
	         : (byte_in == 8'ha9)? 32'hed570001
	         : (byte_in == 8'haa)? 32'he5e80000
	         : (byte_in == 8'hab)? 32'h25a60001
	         : (byte_in == 8'hac)? 32'ha53a0002
	         : (byte_in == 8'had)? 32'h65740003
	         : (byte_in == 8'hae)? 32'h6dcb0002
	         : (byte_in == 8'haf)? 32'had850003
	         : (byte_in == 8'hb0)? 32'hacbd0004
	         : (byte_in == 8'hb1)? 32'h6cf30005
	         : (byte_in == 8'hb2)? 32'h644c0004
	         : (byte_in == 8'hb3)? 32'ha4020005
	         : (byte_in == 8'hb4)? 32'h249e0006
	         : (byte_in == 8'hb5)? 32'he4d00007
	         : (byte_in == 8'hb6)? 32'hec6f0006
	         : (byte_in == 8'hb7)? 32'h2c210007
	         : (byte_in == 8'hb8)? 32'hfd110004
	         : (byte_in == 8'hb9)? 32'h3d5f0005
	         : (byte_in == 8'hba)? 32'h35e00004
	         : (byte_in == 8'hbb)? 32'hf5ae0005
	         : (byte_in == 8'hbc)? 32'h75320006
	         : (byte_in == 8'hbd)? 32'hb57c0007
	         : (byte_in == 8'hbe)? 32'hbdc30006
	         : (byte_in == 8'hbf)? 32'h7d8d0007
	         : (byte_in == 8'hc0)? 32'hbfb20008
	         : (byte_in == 8'hc1)? 32'h7ffc0009
	         : (byte_in == 8'hc2)? 32'h77430008
	         : (byte_in == 8'hc3)? 32'hb70d0009
	         : (byte_in == 8'hc4)? 32'h3791000a
	         : (byte_in == 8'hc5)? 32'hf7df000b
	         : (byte_in == 8'hc6)? 32'hff60000a
	         : (byte_in == 8'hc7)? 32'h3f2e000b
	         : (byte_in == 8'hc8)? 32'hee1e0008
	         : (byte_in == 8'hc9)? 32'h2e500009
	         : (byte_in == 8'hca)? 32'h26ef0008
	         : (byte_in == 8'hcb)? 32'he6a10009
	         : (byte_in == 8'hcc)? 32'h663d000a
	         : (byte_in == 8'hcd)? 32'ha673000b
	         : (byte_in == 8'hce)? 32'haecc000a
	         : (byte_in == 8'hcf)? 32'h6e82000b
	         : (byte_in == 8'hd0)? 32'h6fba000c
	         : (byte_in == 8'hd1)? 32'haff4000d
	         : (byte_in == 8'hd2)? 32'ha74b000c
	         : (byte_in == 8'hd3)? 32'h6705000d
	         : (byte_in == 8'hd4)? 32'he799000e
	         : (byte_in == 8'hd5)? 32'h27d7000f
	         : (byte_in == 8'hd6)? 32'h2f68000e
	         : (byte_in == 8'hd7)? 32'hef26000f
	         : (byte_in == 8'hd8)? 32'h3e16000c
	         : (byte_in == 8'hd9)? 32'hfe58000d
	         : (byte_in == 8'hda)? 32'hf6e7000c
	         : (byte_in == 8'hdb)? 32'h36a9000d
	         : (byte_in == 8'hdc)? 32'hb635000e
	         : (byte_in == 8'hdd)? 32'h767b000f
	         : (byte_in == 8'hde)? 32'h7ec4000e
	         : (byte_in == 8'hdf)? 32'hbe8a000f
	         : (byte_in == 8'he0)? 32'hd41b0008
	         : (byte_in == 8'he1)? 32'h14550009
	         : (byte_in == 8'he2)? 32'h1cea0008
	         : (byte_in == 8'he3)? 32'hdca40009
	         : (byte_in == 8'he4)? 32'h5c38000a
	         : (byte_in == 8'he5)? 32'h9c76000b
	         : (byte_in == 8'he6)? 32'h94c9000a
	         : (byte_in == 8'he7)? 32'h5487000b
	         : (byte_in == 8'he8)? 32'h85b70008
	         : (byte_in == 8'he9)? 32'h45f90009
	         : (byte_in == 8'hea)? 32'h4d460008
	         : (byte_in == 8'heb)? 32'h8d080009
	         : (byte_in == 8'hec)? 32'h0d94000a
	         : (byte_in == 8'hed)? 32'hcdda000b
	         : (byte_in == 8'hee)? 32'hc565000a
	         : (byte_in == 8'hef)? 32'h052b000b
	         : (byte_in == 8'hf0)? 32'h0413000c
	         : (byte_in == 8'hf1)? 32'hc45d000d
	         : (byte_in == 8'hf2)? 32'hcce2000c
	         : (byte_in == 8'hf3)? 32'h0cac000d
	         : (byte_in == 8'hf4)? 32'h8c30000e
	         : (byte_in == 8'hf5)? 32'h4c7e000f
	         : (byte_in == 8'hf6)? 32'h44c1000e
	         : (byte_in == 8'hf7)? 32'h848f000f
	         : (byte_in == 8'hf8)? 32'h55bf000c
	         : (byte_in == 8'hf9)? 32'h95f1000d
	         : (byte_in == 8'hfa)? 32'h9d4e000c
	         : (byte_in == 8'hfb)? 32'h5d00000d
	         : (byte_in == 8'hfc)? 32'hdd9c000e
	         : (byte_in == 8'hfd)? 32'h1dd2000f
	         : (byte_in == 8'hfe)? 32'h156d000e
	         :                     32'hd523000f;

endmodule
//}}}

module TABLE1(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h515c0010
	         : (byte_in == 8'h02)? 32'h2e390000
	         : (byte_in == 8'h03)? 32'h7f650010
	         : (byte_in == 8'h04)? 32'ha2b80020
	         : (byte_in == 8'h05)? 32'hf3e40030
	         : (byte_in == 8'h06)? 32'h8c810020
	         : (byte_in == 8'h07)? 32'hdddd0030
	         : (byte_in == 8'h08)? 32'h5c720000
	         : (byte_in == 8'h09)? 32'h0d2e0010
	         : (byte_in == 8'h0a)? 32'h724b0000
	         : (byte_in == 8'h0b)? 32'h23170010
	         : (byte_in == 8'h0c)? 32'hfeca0020
	         : (byte_in == 8'h0d)? 32'haf960030
	         : (byte_in == 8'h0e)? 32'hd0f30020
	         : (byte_in == 8'h0f)? 32'h81af0030
	         : (byte_in == 8'h10)? 32'h4dce0040
	         : (byte_in == 8'h11)? 32'h1c920050
	         : (byte_in == 8'h12)? 32'h63f70040
	         : (byte_in == 8'h13)? 32'h32ab0050
	         : (byte_in == 8'h14)? 32'hef760060
	         : (byte_in == 8'h15)? 32'hbe2a0070
	         : (byte_in == 8'h16)? 32'hc14f0060
	         : (byte_in == 8'h17)? 32'h90130070
	         : (byte_in == 8'h18)? 32'h11bc0040
	         : (byte_in == 8'h19)? 32'h40e00050
	         : (byte_in == 8'h1a)? 32'h3f850040
	         : (byte_in == 8'h1b)? 32'h6ed90050
	         : (byte_in == 8'h1c)? 32'hb3040060
	         : (byte_in == 8'h1d)? 32'he2580070
	         : (byte_in == 8'h1e)? 32'h9d3d0060
	         : (byte_in == 8'h1f)? 32'hcc610070
	         : (byte_in == 8'h20)? 32'h78ab0000
	         : (byte_in == 8'h21)? 32'h29f70010
	         : (byte_in == 8'h22)? 32'h56920000
	         : (byte_in == 8'h23)? 32'h07ce0010
	         : (byte_in == 8'h24)? 32'hda130020
	         : (byte_in == 8'h25)? 32'h8b4f0030
	         : (byte_in == 8'h26)? 32'hf42a0020
	         : (byte_in == 8'h27)? 32'ha5760030
	         : (byte_in == 8'h28)? 32'h24d90000
	         : (byte_in == 8'h29)? 32'h75850010
	         : (byte_in == 8'h2a)? 32'h0ae00000
	         : (byte_in == 8'h2b)? 32'h5bbc0010
	         : (byte_in == 8'h2c)? 32'h86610020
	         : (byte_in == 8'h2d)? 32'hd73d0030
	         : (byte_in == 8'h2e)? 32'ha8580020
	         : (byte_in == 8'h2f)? 32'hf9040030
	         : (byte_in == 8'h30)? 32'h35650040
	         : (byte_in == 8'h31)? 32'h64390050
	         : (byte_in == 8'h32)? 32'h1b5c0040
	         : (byte_in == 8'h33)? 32'h4a000050
	         : (byte_in == 8'h34)? 32'h97dd0060
	         : (byte_in == 8'h35)? 32'hc6810070
	         : (byte_in == 8'h36)? 32'hb9e40060
	         : (byte_in == 8'h37)? 32'he8b80070
	         : (byte_in == 8'h38)? 32'h69170040
	         : (byte_in == 8'h39)? 32'h384b0050
	         : (byte_in == 8'h3a)? 32'h472e0040
	         : (byte_in == 8'h3b)? 32'h16720050
	         : (byte_in == 8'h3c)? 32'hcbaf0060
	         : (byte_in == 8'h3d)? 32'h9af30070
	         : (byte_in == 8'h3e)? 32'he5960060
	         : (byte_in == 8'h3f)? 32'hb4ca0070
	         : (byte_in == 8'h40)? 32'h5bd20080
	         : (byte_in == 8'h41)? 32'h0a8e0090
	         : (byte_in == 8'h42)? 32'h75eb0080
	         : (byte_in == 8'h43)? 32'h24b70090
	         : (byte_in == 8'h44)? 32'hf96a00a0
	         : (byte_in == 8'h45)? 32'ha83600b0
	         : (byte_in == 8'h46)? 32'hd75300a0
	         : (byte_in == 8'h47)? 32'h860f00b0
	         : (byte_in == 8'h48)? 32'h07a00080
	         : (byte_in == 8'h49)? 32'h56fc0090
	         : (byte_in == 8'h4a)? 32'h29990080
	         : (byte_in == 8'h4b)? 32'h78c50090
	         : (byte_in == 8'h4c)? 32'ha51800a0
	         : (byte_in == 8'h4d)? 32'hf44400b0
	         : (byte_in == 8'h4e)? 32'h8b2100a0
	         : (byte_in == 8'h4f)? 32'hda7d00b0
	         : (byte_in == 8'h50)? 32'h161c00c0
	         : (byte_in == 8'h51)? 32'h474000d0
	         : (byte_in == 8'h52)? 32'h382500c0
	         : (byte_in == 8'h53)? 32'h697900d0
	         : (byte_in == 8'h54)? 32'hb4a400e0
	         : (byte_in == 8'h55)? 32'he5f800f0
	         : (byte_in == 8'h56)? 32'h9a9d00e0
	         : (byte_in == 8'h57)? 32'hcbc100f0
	         : (byte_in == 8'h58)? 32'h4a6e00c0
	         : (byte_in == 8'h59)? 32'h1b3200d0
	         : (byte_in == 8'h5a)? 32'h645700c0
	         : (byte_in == 8'h5b)? 32'h350b00d0
	         : (byte_in == 8'h5c)? 32'he8d600e0
	         : (byte_in == 8'h5d)? 32'hb98a00f0
	         : (byte_in == 8'h5e)? 32'hc6ef00e0
	         : (byte_in == 8'h5f)? 32'h97b300f0
	         : (byte_in == 8'h60)? 32'h23790080
	         : (byte_in == 8'h61)? 32'h72250090
	         : (byte_in == 8'h62)? 32'h0d400080
	         : (byte_in == 8'h63)? 32'h5c1c0090
	         : (byte_in == 8'h64)? 32'h81c100a0
	         : (byte_in == 8'h65)? 32'hd09d00b0
	         : (byte_in == 8'h66)? 32'haff800a0
	         : (byte_in == 8'h67)? 32'hfea400b0
	         : (byte_in == 8'h68)? 32'h7f0b0080
	         : (byte_in == 8'h69)? 32'h2e570090
	         : (byte_in == 8'h6a)? 32'h51320080
	         : (byte_in == 8'h6b)? 32'h006e0090
	         : (byte_in == 8'h6c)? 32'hddb300a0
	         : (byte_in == 8'h6d)? 32'h8cef00b0
	         : (byte_in == 8'h6e)? 32'hf38a00a0
	         : (byte_in == 8'h6f)? 32'ha2d600b0
	         : (byte_in == 8'h70)? 32'h6eb700c0
	         : (byte_in == 8'h71)? 32'h3feb00d0
	         : (byte_in == 8'h72)? 32'h408e00c0
	         : (byte_in == 8'h73)? 32'h11d200d0
	         : (byte_in == 8'h74)? 32'hcc0f00e0
	         : (byte_in == 8'h75)? 32'h9d5300f0
	         : (byte_in == 8'h76)? 32'he23600e0
	         : (byte_in == 8'h77)? 32'hb36a00f0
	         : (byte_in == 8'h78)? 32'h32c500c0
	         : (byte_in == 8'h79)? 32'h639900d0
	         : (byte_in == 8'h7a)? 32'h1cfc00c0
	         : (byte_in == 8'h7b)? 32'h4da000d0
	         : (byte_in == 8'h7c)? 32'h907d00e0
	         : (byte_in == 8'h7d)? 32'hc12100f0
	         : (byte_in == 8'h7e)? 32'hbe4400e0
	         : (byte_in == 8'h7f)? 32'hef1800f0
	         : (byte_in == 8'h80)? 32'h39a60000
	         : (byte_in == 8'h81)? 32'h68fa0010
	         : (byte_in == 8'h82)? 32'h179f0000
	         : (byte_in == 8'h83)? 32'h46c30010
	         : (byte_in == 8'h84)? 32'h9b1e0020
	         : (byte_in == 8'h85)? 32'hca420030
	         : (byte_in == 8'h86)? 32'hb5270020
	         : (byte_in == 8'h87)? 32'he47b0030
	         : (byte_in == 8'h88)? 32'h65d40000
	         : (byte_in == 8'h89)? 32'h34880010
	         : (byte_in == 8'h8a)? 32'h4bed0000
	         : (byte_in == 8'h8b)? 32'h1ab10010
	         : (byte_in == 8'h8c)? 32'hc76c0020
	         : (byte_in == 8'h8d)? 32'h96300030
	         : (byte_in == 8'h8e)? 32'he9550020
	         : (byte_in == 8'h8f)? 32'hb8090030
	         : (byte_in == 8'h90)? 32'h74680040
	         : (byte_in == 8'h91)? 32'h25340050
	         : (byte_in == 8'h92)? 32'h5a510040
	         : (byte_in == 8'h93)? 32'h0b0d0050
	         : (byte_in == 8'h94)? 32'hd6d00060
	         : (byte_in == 8'h95)? 32'h878c0070
	         : (byte_in == 8'h96)? 32'hf8e90060
	         : (byte_in == 8'h97)? 32'ha9b50070
	         : (byte_in == 8'h98)? 32'h281a0040
	         : (byte_in == 8'h99)? 32'h79460050
	         : (byte_in == 8'h9a)? 32'h06230040
	         : (byte_in == 8'h9b)? 32'h577f0050
	         : (byte_in == 8'h9c)? 32'h8aa20060
	         : (byte_in == 8'h9d)? 32'hdbfe0070
	         : (byte_in == 8'h9e)? 32'ha49b0060
	         : (byte_in == 8'h9f)? 32'hf5c70070
	         : (byte_in == 8'ha0)? 32'h410d0000
	         : (byte_in == 8'ha1)? 32'h10510010
	         : (byte_in == 8'ha2)? 32'h6f340000
	         : (byte_in == 8'ha3)? 32'h3e680010
	         : (byte_in == 8'ha4)? 32'he3b50020
	         : (byte_in == 8'ha5)? 32'hb2e90030
	         : (byte_in == 8'ha6)? 32'hcd8c0020
	         : (byte_in == 8'ha7)? 32'h9cd00030
	         : (byte_in == 8'ha8)? 32'h1d7f0000
	         : (byte_in == 8'ha9)? 32'h4c230010
	         : (byte_in == 8'haa)? 32'h33460000
	         : (byte_in == 8'hab)? 32'h621a0010
	         : (byte_in == 8'hac)? 32'hbfc70020
	         : (byte_in == 8'had)? 32'hee9b0030
	         : (byte_in == 8'hae)? 32'h91fe0020
	         : (byte_in == 8'haf)? 32'hc0a20030
	         : (byte_in == 8'hb0)? 32'h0cc30040
	         : (byte_in == 8'hb1)? 32'h5d9f0050
	         : (byte_in == 8'hb2)? 32'h22fa0040
	         : (byte_in == 8'hb3)? 32'h73a60050
	         : (byte_in == 8'hb4)? 32'hae7b0060
	         : (byte_in == 8'hb5)? 32'hff270070
	         : (byte_in == 8'hb6)? 32'h80420060
	         : (byte_in == 8'hb7)? 32'hd11e0070
	         : (byte_in == 8'hb8)? 32'h50b10040
	         : (byte_in == 8'hb9)? 32'h01ed0050
	         : (byte_in == 8'hba)? 32'h7e880040
	         : (byte_in == 8'hbb)? 32'h2fd40050
	         : (byte_in == 8'hbc)? 32'hf2090060
	         : (byte_in == 8'hbd)? 32'ha3550070
	         : (byte_in == 8'hbe)? 32'hdc300060
	         : (byte_in == 8'hbf)? 32'h8d6c0070
	         : (byte_in == 8'hc0)? 32'h62740080
	         : (byte_in == 8'hc1)? 32'h33280090
	         : (byte_in == 8'hc2)? 32'h4c4d0080
	         : (byte_in == 8'hc3)? 32'h1d110090
	         : (byte_in == 8'hc4)? 32'hc0cc00a0
	         : (byte_in == 8'hc5)? 32'h919000b0
	         : (byte_in == 8'hc6)? 32'heef500a0
	         : (byte_in == 8'hc7)? 32'hbfa900b0
	         : (byte_in == 8'hc8)? 32'h3e060080
	         : (byte_in == 8'hc9)? 32'h6f5a0090
	         : (byte_in == 8'hca)? 32'h103f0080
	         : (byte_in == 8'hcb)? 32'h41630090
	         : (byte_in == 8'hcc)? 32'h9cbe00a0
	         : (byte_in == 8'hcd)? 32'hcde200b0
	         : (byte_in == 8'hce)? 32'hb28700a0
	         : (byte_in == 8'hcf)? 32'he3db00b0
	         : (byte_in == 8'hd0)? 32'h2fba00c0
	         : (byte_in == 8'hd1)? 32'h7ee600d0
	         : (byte_in == 8'hd2)? 32'h018300c0
	         : (byte_in == 8'hd3)? 32'h50df00d0
	         : (byte_in == 8'hd4)? 32'h8d0200e0
	         : (byte_in == 8'hd5)? 32'hdc5e00f0
	         : (byte_in == 8'hd6)? 32'ha33b00e0
	         : (byte_in == 8'hd7)? 32'hf26700f0
	         : (byte_in == 8'hd8)? 32'h73c800c0
	         : (byte_in == 8'hd9)? 32'h229400d0
	         : (byte_in == 8'hda)? 32'h5df100c0
	         : (byte_in == 8'hdb)? 32'h0cad00d0
	         : (byte_in == 8'hdc)? 32'hd17000e0
	         : (byte_in == 8'hdd)? 32'h802c00f0
	         : (byte_in == 8'hde)? 32'hff4900e0
	         : (byte_in == 8'hdf)? 32'hae1500f0
	         : (byte_in == 8'he0)? 32'h1adf0080
	         : (byte_in == 8'he1)? 32'h4b830090
	         : (byte_in == 8'he2)? 32'h34e60080
	         : (byte_in == 8'he3)? 32'h65ba0090
	         : (byte_in == 8'he4)? 32'hb86700a0
	         : (byte_in == 8'he5)? 32'he93b00b0
	         : (byte_in == 8'he6)? 32'h965e00a0
	         : (byte_in == 8'he7)? 32'hc70200b0
	         : (byte_in == 8'he8)? 32'h46ad0080
	         : (byte_in == 8'he9)? 32'h17f10090
	         : (byte_in == 8'hea)? 32'h68940080
	         : (byte_in == 8'heb)? 32'h39c80090
	         : (byte_in == 8'hec)? 32'he41500a0
	         : (byte_in == 8'hed)? 32'hb54900b0
	         : (byte_in == 8'hee)? 32'hca2c00a0
	         : (byte_in == 8'hef)? 32'h9b7000b0
	         : (byte_in == 8'hf0)? 32'h571100c0
	         : (byte_in == 8'hf1)? 32'h064d00d0
	         : (byte_in == 8'hf2)? 32'h792800c0
	         : (byte_in == 8'hf3)? 32'h287400d0
	         : (byte_in == 8'hf4)? 32'hf5a900e0
	         : (byte_in == 8'hf5)? 32'ha4f500f0
	         : (byte_in == 8'hf6)? 32'hdb9000e0
	         : (byte_in == 8'hf7)? 32'h8acc00f0
	         : (byte_in == 8'hf8)? 32'h0b6300c0
	         : (byte_in == 8'hf9)? 32'h5a3f00d0
	         : (byte_in == 8'hfa)? 32'h255a00c0
	         : (byte_in == 8'hfb)? 32'h740600d0
	         : (byte_in == 8'hfc)? 32'ha9db00e0
	         : (byte_in == 8'hfd)? 32'hf88700f0
	         : (byte_in == 8'hfe)? 32'h87e200e0
	         :                     32'hd6be00f0;

endmodule
//}}}

module TABLE2(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'hb7a40100
	         : (byte_in == 8'h02)? 32'h734c0000
	         : (byte_in == 8'h03)? 32'hc4e80100
	         : (byte_in == 8'h04)? 32'ha7b80200
	         : (byte_in == 8'h05)? 32'h101c0300
	         : (byte_in == 8'h06)? 32'hd4f40200
	         : (byte_in == 8'h07)? 32'h63500300
	         : (byte_in == 8'h08)? 32'hee260000
	         : (byte_in == 8'h09)? 32'h59820100
	         : (byte_in == 8'h0a)? 32'h9d6a0000
	         : (byte_in == 8'h0b)? 32'h2ace0100
	         : (byte_in == 8'h0c)? 32'h499e0200
	         : (byte_in == 8'h0d)? 32'hfe3a0300
	         : (byte_in == 8'h0e)? 32'h3ad20200
	         : (byte_in == 8'h0f)? 32'h8d760300
	         : (byte_in == 8'h10)? 32'h8f3e0400
	         : (byte_in == 8'h11)? 32'h389a0500
	         : (byte_in == 8'h12)? 32'hfc720400
	         : (byte_in == 8'h13)? 32'h4bd60500
	         : (byte_in == 8'h14)? 32'h28860600
	         : (byte_in == 8'h15)? 32'h9f220700
	         : (byte_in == 8'h16)? 32'h5bca0600
	         : (byte_in == 8'h17)? 32'hec6e0700
	         : (byte_in == 8'h18)? 32'h61180400
	         : (byte_in == 8'h19)? 32'hd6bc0500
	         : (byte_in == 8'h1a)? 32'h12540400
	         : (byte_in == 8'h1b)? 32'ha5f00500
	         : (byte_in == 8'h1c)? 32'hc6a00600
	         : (byte_in == 8'h1d)? 32'h71040700
	         : (byte_in == 8'h1e)? 32'hb5ec0600
	         : (byte_in == 8'h1f)? 32'h02480700
	         : (byte_in == 8'h20)? 32'h14bd0000
	         : (byte_in == 8'h21)? 32'ha3190100
	         : (byte_in == 8'h22)? 32'h67f10000
	         : (byte_in == 8'h23)? 32'hd0550100
	         : (byte_in == 8'h24)? 32'hb3050200
	         : (byte_in == 8'h25)? 32'h04a10300
	         : (byte_in == 8'h26)? 32'hc0490200
	         : (byte_in == 8'h27)? 32'h77ed0300
	         : (byte_in == 8'h28)? 32'hfa9b0000
	         : (byte_in == 8'h29)? 32'h4d3f0100
	         : (byte_in == 8'h2a)? 32'h89d70000
	         : (byte_in == 8'h2b)? 32'h3e730100
	         : (byte_in == 8'h2c)? 32'h5d230200
	         : (byte_in == 8'h2d)? 32'hea870300
	         : (byte_in == 8'h2e)? 32'h2e6f0200
	         : (byte_in == 8'h2f)? 32'h99cb0300
	         : (byte_in == 8'h30)? 32'h9b830400
	         : (byte_in == 8'h31)? 32'h2c270500
	         : (byte_in == 8'h32)? 32'he8cf0400
	         : (byte_in == 8'h33)? 32'h5f6b0500
	         : (byte_in == 8'h34)? 32'h3c3b0600
	         : (byte_in == 8'h35)? 32'h8b9f0700
	         : (byte_in == 8'h36)? 32'h4f770600
	         : (byte_in == 8'h37)? 32'hf8d30700
	         : (byte_in == 8'h38)? 32'h75a50400
	         : (byte_in == 8'h39)? 32'hc2010500
	         : (byte_in == 8'h3a)? 32'h06e90400
	         : (byte_in == 8'h3b)? 32'hb14d0500
	         : (byte_in == 8'h3c)? 32'hd21d0600
	         : (byte_in == 8'h3d)? 32'h65b90700
	         : (byte_in == 8'h3e)? 32'ha1510600
	         : (byte_in == 8'h3f)? 32'h16f50700
	         : (byte_in == 8'h40)? 32'hde320800
	         : (byte_in == 8'h41)? 32'h69960900
	         : (byte_in == 8'h42)? 32'had7e0800
	         : (byte_in == 8'h43)? 32'h1ada0900
	         : (byte_in == 8'h44)? 32'h798a0a00
	         : (byte_in == 8'h45)? 32'hce2e0b00
	         : (byte_in == 8'h46)? 32'h0ac60a00
	         : (byte_in == 8'h47)? 32'hbd620b00
	         : (byte_in == 8'h48)? 32'h30140800
	         : (byte_in == 8'h49)? 32'h87b00900
	         : (byte_in == 8'h4a)? 32'h43580800
	         : (byte_in == 8'h4b)? 32'hf4fc0900
	         : (byte_in == 8'h4c)? 32'h97ac0a00
	         : (byte_in == 8'h4d)? 32'h20080b00
	         : (byte_in == 8'h4e)? 32'he4e00a00
	         : (byte_in == 8'h4f)? 32'h53440b00
	         : (byte_in == 8'h50)? 32'h510c0c00
	         : (byte_in == 8'h51)? 32'he6a80d00
	         : (byte_in == 8'h52)? 32'h22400c00
	         : (byte_in == 8'h53)? 32'h95e40d00
	         : (byte_in == 8'h54)? 32'hf6b40e00
	         : (byte_in == 8'h55)? 32'h41100f00
	         : (byte_in == 8'h56)? 32'h85f80e00
	         : (byte_in == 8'h57)? 32'h325c0f00
	         : (byte_in == 8'h58)? 32'hbf2a0c00
	         : (byte_in == 8'h59)? 32'h088e0d00
	         : (byte_in == 8'h5a)? 32'hcc660c00
	         : (byte_in == 8'h5b)? 32'h7bc20d00
	         : (byte_in == 8'h5c)? 32'h18920e00
	         : (byte_in == 8'h5d)? 32'haf360f00
	         : (byte_in == 8'h5e)? 32'h6bde0e00
	         : (byte_in == 8'h5f)? 32'hdc7a0f00
	         : (byte_in == 8'h60)? 32'hca8f0800
	         : (byte_in == 8'h61)? 32'h7d2b0900
	         : (byte_in == 8'h62)? 32'hb9c30800
	         : (byte_in == 8'h63)? 32'h0e670900
	         : (byte_in == 8'h64)? 32'h6d370a00
	         : (byte_in == 8'h65)? 32'hda930b00
	         : (byte_in == 8'h66)? 32'h1e7b0a00
	         : (byte_in == 8'h67)? 32'ha9df0b00
	         : (byte_in == 8'h68)? 32'h24a90800
	         : (byte_in == 8'h69)? 32'h930d0900
	         : (byte_in == 8'h6a)? 32'h57e50800
	         : (byte_in == 8'h6b)? 32'he0410900
	         : (byte_in == 8'h6c)? 32'h83110a00
	         : (byte_in == 8'h6d)? 32'h34b50b00
	         : (byte_in == 8'h6e)? 32'hf05d0a00
	         : (byte_in == 8'h6f)? 32'h47f90b00
	         : (byte_in == 8'h70)? 32'h45b10c00
	         : (byte_in == 8'h71)? 32'hf2150d00
	         : (byte_in == 8'h72)? 32'h36fd0c00
	         : (byte_in == 8'h73)? 32'h81590d00
	         : (byte_in == 8'h74)? 32'he2090e00
	         : (byte_in == 8'h75)? 32'h55ad0f00
	         : (byte_in == 8'h76)? 32'h91450e00
	         : (byte_in == 8'h77)? 32'h26e10f00
	         : (byte_in == 8'h78)? 32'hab970c00
	         : (byte_in == 8'h79)? 32'h1c330d00
	         : (byte_in == 8'h7a)? 32'hd8db0c00
	         : (byte_in == 8'h7b)? 32'h6f7f0d00
	         : (byte_in == 8'h7c)? 32'h0c2f0e00
	         : (byte_in == 8'h7d)? 32'hbb8b0f00
	         : (byte_in == 8'h7e)? 32'h7f630e00
	         : (byte_in == 8'h7f)? 32'hc8c70f00
	         : (byte_in == 8'h80)? 32'he18b0000
	         : (byte_in == 8'h81)? 32'h562f0100
	         : (byte_in == 8'h82)? 32'h92c70000
	         : (byte_in == 8'h83)? 32'h25630100
	         : (byte_in == 8'h84)? 32'h46330200
	         : (byte_in == 8'h85)? 32'hf1970300
	         : (byte_in == 8'h86)? 32'h357f0200
	         : (byte_in == 8'h87)? 32'h82db0300
	         : (byte_in == 8'h88)? 32'h0fad0000
	         : (byte_in == 8'h89)? 32'hb8090100
	         : (byte_in == 8'h8a)? 32'h7ce10000
	         : (byte_in == 8'h8b)? 32'hcb450100
	         : (byte_in == 8'h8c)? 32'ha8150200
	         : (byte_in == 8'h8d)? 32'h1fb10300
	         : (byte_in == 8'h8e)? 32'hdb590200
	         : (byte_in == 8'h8f)? 32'h6cfd0300
	         : (byte_in == 8'h90)? 32'h6eb50400
	         : (byte_in == 8'h91)? 32'hd9110500
	         : (byte_in == 8'h92)? 32'h1df90400
	         : (byte_in == 8'h93)? 32'haa5d0500
	         : (byte_in == 8'h94)? 32'hc90d0600
	         : (byte_in == 8'h95)? 32'h7ea90700
	         : (byte_in == 8'h96)? 32'hba410600
	         : (byte_in == 8'h97)? 32'h0de50700
	         : (byte_in == 8'h98)? 32'h80930400
	         : (byte_in == 8'h99)? 32'h37370500
	         : (byte_in == 8'h9a)? 32'hf3df0400
	         : (byte_in == 8'h9b)? 32'h447b0500
	         : (byte_in == 8'h9c)? 32'h272b0600
	         : (byte_in == 8'h9d)? 32'h908f0700
	         : (byte_in == 8'h9e)? 32'h54670600
	         : (byte_in == 8'h9f)? 32'he3c30700
	         : (byte_in == 8'ha0)? 32'hf5360000
	         : (byte_in == 8'ha1)? 32'h42920100
	         : (byte_in == 8'ha2)? 32'h867a0000
	         : (byte_in == 8'ha3)? 32'h31de0100
	         : (byte_in == 8'ha4)? 32'h528e0200
	         : (byte_in == 8'ha5)? 32'he52a0300
	         : (byte_in == 8'ha6)? 32'h21c20200
	         : (byte_in == 8'ha7)? 32'h96660300
	         : (byte_in == 8'ha8)? 32'h1b100000
	         : (byte_in == 8'ha9)? 32'hacb40100
	         : (byte_in == 8'haa)? 32'h685c0000
	         : (byte_in == 8'hab)? 32'hdff80100
	         : (byte_in == 8'hac)? 32'hbca80200
	         : (byte_in == 8'had)? 32'h0b0c0300
	         : (byte_in == 8'hae)? 32'hcfe40200
	         : (byte_in == 8'haf)? 32'h78400300
	         : (byte_in == 8'hb0)? 32'h7a080400
	         : (byte_in == 8'hb1)? 32'hcdac0500
	         : (byte_in == 8'hb2)? 32'h09440400
	         : (byte_in == 8'hb3)? 32'hbee00500
	         : (byte_in == 8'hb4)? 32'hddb00600
	         : (byte_in == 8'hb5)? 32'h6a140700
	         : (byte_in == 8'hb6)? 32'haefc0600
	         : (byte_in == 8'hb7)? 32'h19580700
	         : (byte_in == 8'hb8)? 32'h942e0400
	         : (byte_in == 8'hb9)? 32'h238a0500
	         : (byte_in == 8'hba)? 32'he7620400
	         : (byte_in == 8'hbb)? 32'h50c60500
	         : (byte_in == 8'hbc)? 32'h33960600
	         : (byte_in == 8'hbd)? 32'h84320700
	         : (byte_in == 8'hbe)? 32'h40da0600
	         : (byte_in == 8'hbf)? 32'hf77e0700
	         : (byte_in == 8'hc0)? 32'h3fb90800
	         : (byte_in == 8'hc1)? 32'h881d0900
	         : (byte_in == 8'hc2)? 32'h4cf50800
	         : (byte_in == 8'hc3)? 32'hfb510900
	         : (byte_in == 8'hc4)? 32'h98010a00
	         : (byte_in == 8'hc5)? 32'h2fa50b00
	         : (byte_in == 8'hc6)? 32'heb4d0a00
	         : (byte_in == 8'hc7)? 32'h5ce90b00
	         : (byte_in == 8'hc8)? 32'hd19f0800
	         : (byte_in == 8'hc9)? 32'h663b0900
	         : (byte_in == 8'hca)? 32'ha2d30800
	         : (byte_in == 8'hcb)? 32'h15770900
	         : (byte_in == 8'hcc)? 32'h76270a00
	         : (byte_in == 8'hcd)? 32'hc1830b00
	         : (byte_in == 8'hce)? 32'h056b0a00
	         : (byte_in == 8'hcf)? 32'hb2cf0b00
	         : (byte_in == 8'hd0)? 32'hb0870c00
	         : (byte_in == 8'hd1)? 32'h07230d00
	         : (byte_in == 8'hd2)? 32'hc3cb0c00
	         : (byte_in == 8'hd3)? 32'h746f0d00
	         : (byte_in == 8'hd4)? 32'h173f0e00
	         : (byte_in == 8'hd5)? 32'ha09b0f00
	         : (byte_in == 8'hd6)? 32'h64730e00
	         : (byte_in == 8'hd7)? 32'hd3d70f00
	         : (byte_in == 8'hd8)? 32'h5ea10c00
	         : (byte_in == 8'hd9)? 32'he9050d00
	         : (byte_in == 8'hda)? 32'h2ded0c00
	         : (byte_in == 8'hdb)? 32'h9a490d00
	         : (byte_in == 8'hdc)? 32'hf9190e00
	         : (byte_in == 8'hdd)? 32'h4ebd0f00
	         : (byte_in == 8'hde)? 32'h8a550e00
	         : (byte_in == 8'hdf)? 32'h3df10f00
	         : (byte_in == 8'he0)? 32'h2b040800
	         : (byte_in == 8'he1)? 32'h9ca00900
	         : (byte_in == 8'he2)? 32'h58480800
	         : (byte_in == 8'he3)? 32'hefec0900
	         : (byte_in == 8'he4)? 32'h8cbc0a00
	         : (byte_in == 8'he5)? 32'h3b180b00
	         : (byte_in == 8'he6)? 32'hfff00a00
	         : (byte_in == 8'he7)? 32'h48540b00
	         : (byte_in == 8'he8)? 32'hc5220800
	         : (byte_in == 8'he9)? 32'h72860900
	         : (byte_in == 8'hea)? 32'hb66e0800
	         : (byte_in == 8'heb)? 32'h01ca0900
	         : (byte_in == 8'hec)? 32'h629a0a00
	         : (byte_in == 8'hed)? 32'hd53e0b00
	         : (byte_in == 8'hee)? 32'h11d60a00
	         : (byte_in == 8'hef)? 32'ha6720b00
	         : (byte_in == 8'hf0)? 32'ha43a0c00
	         : (byte_in == 8'hf1)? 32'h139e0d00
	         : (byte_in == 8'hf2)? 32'hd7760c00
	         : (byte_in == 8'hf3)? 32'h60d20d00
	         : (byte_in == 8'hf4)? 32'h03820e00
	         : (byte_in == 8'hf5)? 32'hb4260f00
	         : (byte_in == 8'hf6)? 32'h70ce0e00
	         : (byte_in == 8'hf7)? 32'hc76a0f00
	         : (byte_in == 8'hf8)? 32'h4a1c0c00
	         : (byte_in == 8'hf9)? 32'hfdb80d00
	         : (byte_in == 8'hfa)? 32'h39500c00
	         : (byte_in == 8'hfb)? 32'h8ef40d00
	         : (byte_in == 8'hfc)? 32'heda40e00
	         : (byte_in == 8'hfd)? 32'h5a000f00
	         : (byte_in == 8'hfe)? 32'h9ee80e00
	         :                     32'h294c0f00;

endmodule
//}}}

module TABLE3(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h74951000
	         : (byte_in == 8'h02)? 32'hcba90000
	         : (byte_in == 8'h03)? 32'hbf3c1000
	         : (byte_in == 8'h04)? 32'he92a2000
	         : (byte_in == 8'h05)? 32'h9dbf3000
	         : (byte_in == 8'h06)? 32'h22832000
	         : (byte_in == 8'h07)? 32'h56163000
	         : (byte_in == 8'h08)? 32'h97530000
	         : (byte_in == 8'h09)? 32'he3c61000
	         : (byte_in == 8'h0a)? 32'h5cfa0000
	         : (byte_in == 8'h0b)? 32'h286f1000
	         : (byte_in == 8'h0c)? 32'h7e792000
	         : (byte_in == 8'h0d)? 32'h0aec3000
	         : (byte_in == 8'h0e)? 32'hb5d02000
	         : (byte_in == 8'h0f)? 32'hc1453000
	         : (byte_in == 8'h10)? 32'h121b4000
	         : (byte_in == 8'h11)? 32'h668e5000
	         : (byte_in == 8'h12)? 32'hd9b24000
	         : (byte_in == 8'h13)? 32'had275000
	         : (byte_in == 8'h14)? 32'hfb316000
	         : (byte_in == 8'h15)? 32'h8fa47000
	         : (byte_in == 8'h16)? 32'h30986000
	         : (byte_in == 8'h17)? 32'h440d7000
	         : (byte_in == 8'h18)? 32'h85484000
	         : (byte_in == 8'h19)? 32'hf1dd5000
	         : (byte_in == 8'h1a)? 32'h4ee14000
	         : (byte_in == 8'h1b)? 32'h3a745000
	         : (byte_in == 8'h1c)? 32'h6c626000
	         : (byte_in == 8'h1d)? 32'h18f77000
	         : (byte_in == 8'h1e)? 32'ha7cb6000
	         : (byte_in == 8'h1f)? 32'hd35e7000
	         : (byte_in == 8'h20)? 32'he6570000
	         : (byte_in == 8'h21)? 32'h92c21000
	         : (byte_in == 8'h22)? 32'h2dfe0000
	         : (byte_in == 8'h23)? 32'h596b1000
	         : (byte_in == 8'h24)? 32'h0f7d2000
	         : (byte_in == 8'h25)? 32'h7be83000
	         : (byte_in == 8'h26)? 32'hc4d42000
	         : (byte_in == 8'h27)? 32'hb0413000
	         : (byte_in == 8'h28)? 32'h71040000
	         : (byte_in == 8'h29)? 32'h05911000
	         : (byte_in == 8'h2a)? 32'hbaad0000
	         : (byte_in == 8'h2b)? 32'hce381000
	         : (byte_in == 8'h2c)? 32'h982e2000
	         : (byte_in == 8'h2d)? 32'hecbb3000
	         : (byte_in == 8'h2e)? 32'h53872000
	         : (byte_in == 8'h2f)? 32'h27123000
	         : (byte_in == 8'h30)? 32'hf44c4000
	         : (byte_in == 8'h31)? 32'h80d95000
	         : (byte_in == 8'h32)? 32'h3fe54000
	         : (byte_in == 8'h33)? 32'h4b705000
	         : (byte_in == 8'h34)? 32'h1d666000
	         : (byte_in == 8'h35)? 32'h69f37000
	         : (byte_in == 8'h36)? 32'hd6cf6000
	         : (byte_in == 8'h37)? 32'ha25a7000
	         : (byte_in == 8'h38)? 32'h631f4000
	         : (byte_in == 8'h39)? 32'h178a5000
	         : (byte_in == 8'h3a)? 32'ha8b64000
	         : (byte_in == 8'h3b)? 32'hdc235000
	         : (byte_in == 8'h3c)? 32'h8a356000
	         : (byte_in == 8'h3d)? 32'hfea07000
	         : (byte_in == 8'h3e)? 32'h419c6000
	         : (byte_in == 8'h3f)? 32'h35097000
	         : (byte_in == 8'h40)? 32'he4788000
	         : (byte_in == 8'h41)? 32'h90ed9000
	         : (byte_in == 8'h42)? 32'h2fd18000
	         : (byte_in == 8'h43)? 32'h5b449000
	         : (byte_in == 8'h44)? 32'h0d52a000
	         : (byte_in == 8'h45)? 32'h79c7b000
	         : (byte_in == 8'h46)? 32'hc6fba000
	         : (byte_in == 8'h47)? 32'hb26eb000
	         : (byte_in == 8'h48)? 32'h732b8000
	         : (byte_in == 8'h49)? 32'h07be9000
	         : (byte_in == 8'h4a)? 32'hb8828000
	         : (byte_in == 8'h4b)? 32'hcc179000
	         : (byte_in == 8'h4c)? 32'h9a01a000
	         : (byte_in == 8'h4d)? 32'hee94b000
	         : (byte_in == 8'h4e)? 32'h51a8a000
	         : (byte_in == 8'h4f)? 32'h253db000
	         : (byte_in == 8'h50)? 32'hf663c000
	         : (byte_in == 8'h51)? 32'h82f6d000
	         : (byte_in == 8'h52)? 32'h3dcac000
	         : (byte_in == 8'h53)? 32'h495fd000
	         : (byte_in == 8'h54)? 32'h1f49e000
	         : (byte_in == 8'h55)? 32'h6bdcf000
	         : (byte_in == 8'h56)? 32'hd4e0e000
	         : (byte_in == 8'h57)? 32'ha075f000
	         : (byte_in == 8'h58)? 32'h6130c000
	         : (byte_in == 8'h59)? 32'h15a5d000
	         : (byte_in == 8'h5a)? 32'haa99c000
	         : (byte_in == 8'h5b)? 32'hde0cd000
	         : (byte_in == 8'h5c)? 32'h881ae000
	         : (byte_in == 8'h5d)? 32'hfc8ff000
	         : (byte_in == 8'h5e)? 32'h43b3e000
	         : (byte_in == 8'h5f)? 32'h3726f000
	         : (byte_in == 8'h60)? 32'h022f8000
	         : (byte_in == 8'h61)? 32'h76ba9000
	         : (byte_in == 8'h62)? 32'hc9868000
	         : (byte_in == 8'h63)? 32'hbd139000
	         : (byte_in == 8'h64)? 32'heb05a000
	         : (byte_in == 8'h65)? 32'h9f90b000
	         : (byte_in == 8'h66)? 32'h20aca000
	         : (byte_in == 8'h67)? 32'h5439b000
	         : (byte_in == 8'h68)? 32'h957c8000
	         : (byte_in == 8'h69)? 32'he1e99000
	         : (byte_in == 8'h6a)? 32'h5ed58000
	         : (byte_in == 8'h6b)? 32'h2a409000
	         : (byte_in == 8'h6c)? 32'h7c56a000
	         : (byte_in == 8'h6d)? 32'h08c3b000
	         : (byte_in == 8'h6e)? 32'hb7ffa000
	         : (byte_in == 8'h6f)? 32'hc36ab000
	         : (byte_in == 8'h70)? 32'h1034c000
	         : (byte_in == 8'h71)? 32'h64a1d000
	         : (byte_in == 8'h72)? 32'hdb9dc000
	         : (byte_in == 8'h73)? 32'haf08d000
	         : (byte_in == 8'h74)? 32'hf91ee000
	         : (byte_in == 8'h75)? 32'h8d8bf000
	         : (byte_in == 8'h76)? 32'h32b7e000
	         : (byte_in == 8'h77)? 32'h4622f000
	         : (byte_in == 8'h78)? 32'h8767c000
	         : (byte_in == 8'h79)? 32'hf3f2d000
	         : (byte_in == 8'h7a)? 32'h4ccec000
	         : (byte_in == 8'h7b)? 32'h385bd000
	         : (byte_in == 8'h7c)? 32'h6e4de000
	         : (byte_in == 8'h7d)? 32'h1ad8f000
	         : (byte_in == 8'h7e)? 32'ha5e4e000
	         : (byte_in == 8'h7f)? 32'hd171f000
	         : (byte_in == 8'h80)? 32'h045f0000
	         : (byte_in == 8'h81)? 32'h70ca1000
	         : (byte_in == 8'h82)? 32'hcff60000
	         : (byte_in == 8'h83)? 32'hbb631000
	         : (byte_in == 8'h84)? 32'hed752000
	         : (byte_in == 8'h85)? 32'h99e03000
	         : (byte_in == 8'h86)? 32'h26dc2000
	         : (byte_in == 8'h87)? 32'h52493000
	         : (byte_in == 8'h88)? 32'h930c0000
	         : (byte_in == 8'h89)? 32'he7991000
	         : (byte_in == 8'h8a)? 32'h58a50000
	         : (byte_in == 8'h8b)? 32'h2c301000
	         : (byte_in == 8'h8c)? 32'h7a262000
	         : (byte_in == 8'h8d)? 32'h0eb33000
	         : (byte_in == 8'h8e)? 32'hb18f2000
	         : (byte_in == 8'h8f)? 32'hc51a3000
	         : (byte_in == 8'h90)? 32'h16444000
	         : (byte_in == 8'h91)? 32'h62d15000
	         : (byte_in == 8'h92)? 32'hdded4000
	         : (byte_in == 8'h93)? 32'ha9785000
	         : (byte_in == 8'h94)? 32'hff6e6000
	         : (byte_in == 8'h95)? 32'h8bfb7000
	         : (byte_in == 8'h96)? 32'h34c76000
	         : (byte_in == 8'h97)? 32'h40527000
	         : (byte_in == 8'h98)? 32'h81174000
	         : (byte_in == 8'h99)? 32'hf5825000
	         : (byte_in == 8'h9a)? 32'h4abe4000
	         : (byte_in == 8'h9b)? 32'h3e2b5000
	         : (byte_in == 8'h9c)? 32'h683d6000
	         : (byte_in == 8'h9d)? 32'h1ca87000
	         : (byte_in == 8'h9e)? 32'ha3946000
	         : (byte_in == 8'h9f)? 32'hd7017000
	         : (byte_in == 8'ha0)? 32'he2080000
	         : (byte_in == 8'ha1)? 32'h969d1000
	         : (byte_in == 8'ha2)? 32'h29a10000
	         : (byte_in == 8'ha3)? 32'h5d341000
	         : (byte_in == 8'ha4)? 32'h0b222000
	         : (byte_in == 8'ha5)? 32'h7fb73000
	         : (byte_in == 8'ha6)? 32'hc08b2000
	         : (byte_in == 8'ha7)? 32'hb41e3000
	         : (byte_in == 8'ha8)? 32'h755b0000
	         : (byte_in == 8'ha9)? 32'h01ce1000
	         : (byte_in == 8'haa)? 32'hbef20000
	         : (byte_in == 8'hab)? 32'hca671000
	         : (byte_in == 8'hac)? 32'h9c712000
	         : (byte_in == 8'had)? 32'he8e43000
	         : (byte_in == 8'hae)? 32'h57d82000
	         : (byte_in == 8'haf)? 32'h234d3000
	         : (byte_in == 8'hb0)? 32'hf0134000
	         : (byte_in == 8'hb1)? 32'h84865000
	         : (byte_in == 8'hb2)? 32'h3bba4000
	         : (byte_in == 8'hb3)? 32'h4f2f5000
	         : (byte_in == 8'hb4)? 32'h19396000
	         : (byte_in == 8'hb5)? 32'h6dac7000
	         : (byte_in == 8'hb6)? 32'hd2906000
	         : (byte_in == 8'hb7)? 32'ha6057000
	         : (byte_in == 8'hb8)? 32'h67404000
	         : (byte_in == 8'hb9)? 32'h13d55000
	         : (byte_in == 8'hba)? 32'hace94000
	         : (byte_in == 8'hbb)? 32'hd87c5000
	         : (byte_in == 8'hbc)? 32'h8e6a6000
	         : (byte_in == 8'hbd)? 32'hfaff7000
	         : (byte_in == 8'hbe)? 32'h45c36000
	         : (byte_in == 8'hbf)? 32'h31567000
	         : (byte_in == 8'hc0)? 32'he0278000
	         : (byte_in == 8'hc1)? 32'h94b29000
	         : (byte_in == 8'hc2)? 32'h2b8e8000
	         : (byte_in == 8'hc3)? 32'h5f1b9000
	         : (byte_in == 8'hc4)? 32'h090da000
	         : (byte_in == 8'hc5)? 32'h7d98b000
	         : (byte_in == 8'hc6)? 32'hc2a4a000
	         : (byte_in == 8'hc7)? 32'hb631b000
	         : (byte_in == 8'hc8)? 32'h77748000
	         : (byte_in == 8'hc9)? 32'h03e19000
	         : (byte_in == 8'hca)? 32'hbcdd8000
	         : (byte_in == 8'hcb)? 32'hc8489000
	         : (byte_in == 8'hcc)? 32'h9e5ea000
	         : (byte_in == 8'hcd)? 32'heacbb000
	         : (byte_in == 8'hce)? 32'h55f7a000
	         : (byte_in == 8'hcf)? 32'h2162b000
	         : (byte_in == 8'hd0)? 32'hf23cc000
	         : (byte_in == 8'hd1)? 32'h86a9d000
	         : (byte_in == 8'hd2)? 32'h3995c000
	         : (byte_in == 8'hd3)? 32'h4d00d000
	         : (byte_in == 8'hd4)? 32'h1b16e000
	         : (byte_in == 8'hd5)? 32'h6f83f000
	         : (byte_in == 8'hd6)? 32'hd0bfe000
	         : (byte_in == 8'hd7)? 32'ha42af000
	         : (byte_in == 8'hd8)? 32'h656fc000
	         : (byte_in == 8'hd9)? 32'h11fad000
	         : (byte_in == 8'hda)? 32'haec6c000
	         : (byte_in == 8'hdb)? 32'hda53d000
	         : (byte_in == 8'hdc)? 32'h8c45e000
	         : (byte_in == 8'hdd)? 32'hf8d0f000
	         : (byte_in == 8'hde)? 32'h47ece000
	         : (byte_in == 8'hdf)? 32'h3379f000
	         : (byte_in == 8'he0)? 32'h06708000
	         : (byte_in == 8'he1)? 32'h72e59000
	         : (byte_in == 8'he2)? 32'hcdd98000
	         : (byte_in == 8'he3)? 32'hb94c9000
	         : (byte_in == 8'he4)? 32'hef5aa000
	         : (byte_in == 8'he5)? 32'h9bcfb000
	         : (byte_in == 8'he6)? 32'h24f3a000
	         : (byte_in == 8'he7)? 32'h5066b000
	         : (byte_in == 8'he8)? 32'h91238000
	         : (byte_in == 8'he9)? 32'he5b69000
	         : (byte_in == 8'hea)? 32'h5a8a8000
	         : (byte_in == 8'heb)? 32'h2e1f9000
	         : (byte_in == 8'hec)? 32'h7809a000
	         : (byte_in == 8'hed)? 32'h0c9cb000
	         : (byte_in == 8'hee)? 32'hb3a0a000
	         : (byte_in == 8'hef)? 32'hc735b000
	         : (byte_in == 8'hf0)? 32'h146bc000
	         : (byte_in == 8'hf1)? 32'h60fed000
	         : (byte_in == 8'hf2)? 32'hdfc2c000
	         : (byte_in == 8'hf3)? 32'hab57d000
	         : (byte_in == 8'hf4)? 32'hfd41e000
	         : (byte_in == 8'hf5)? 32'h89d4f000
	         : (byte_in == 8'hf6)? 32'h36e8e000
	         : (byte_in == 8'hf7)? 32'h427df000
	         : (byte_in == 8'hf8)? 32'h8338c000
	         : (byte_in == 8'hf9)? 32'hf7add000
	         : (byte_in == 8'hfa)? 32'h4891c000
	         : (byte_in == 8'hfb)? 32'h3c04d000
	         : (byte_in == 8'hfc)? 32'h6a12e000
	         : (byte_in == 8'hfd)? 32'h1e87f000
	         : (byte_in == 8'hfe)? 32'ha1bbe000
	         :                     32'hd52ef000;

endmodule
//}}}

module TABLE4(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h33b9c010
	         : (byte_in == 8'h02)? 32'h0b2de782
	         : (byte_in == 8'h03)? 32'h38942792
	         : (byte_in == 8'h04)? 32'h5fe7a7b3
	         : (byte_in == 8'h05)? 32'h6c5e67a3
	         : (byte_in == 8'h06)? 32'h54ca4031
	         : (byte_in == 8'h07)? 32'h67738021
	         : (byte_in == 8'h08)? 32'h25e30f14
	         : (byte_in == 8'h09)? 32'h165acf04
	         : (byte_in == 8'h0a)? 32'h2ecee896
	         : (byte_in == 8'h0b)? 32'h1d772886
	         : (byte_in == 8'h0c)? 32'h7a04a8a7
	         : (byte_in == 8'h0d)? 32'h49bd68b7
	         : (byte_in == 8'h0e)? 32'h71294f25
	         : (byte_in == 8'h0f)? 32'h42908f35
	         : (byte_in == 8'h10)? 32'h8c768f77
	         : (byte_in == 8'h11)? 32'hbfcf4f67
	         : (byte_in == 8'h12)? 32'h875b68f5
	         : (byte_in == 8'h13)? 32'hb4e2a8e5
	         : (byte_in == 8'h14)? 32'hd39128c4
	         : (byte_in == 8'h15)? 32'he028e8d4
	         : (byte_in == 8'h16)? 32'hd8bccf46
	         : (byte_in == 8'h17)? 32'heb050f56
	         : (byte_in == 8'h18)? 32'ha9958063
	         : (byte_in == 8'h19)? 32'h9a2c4073
	         : (byte_in == 8'h1a)? 32'ha2b867e1
	         : (byte_in == 8'h1b)? 32'h9101a7f1
	         : (byte_in == 8'h1c)? 32'hf67227d0
	         : (byte_in == 8'h1d)? 32'hc5cbe7c0
	         : (byte_in == 8'h1e)? 32'hfd5fc052
	         : (byte_in == 8'h1f)? 32'hcee60042
	         : (byte_in == 8'h20)? 32'h40ebf9aa
	         : (byte_in == 8'h21)? 32'h735239ba
	         : (byte_in == 8'h22)? 32'h4bc61e28
	         : (byte_in == 8'h23)? 32'h787fde38
	         : (byte_in == 8'h24)? 32'h1f0c5e19
	         : (byte_in == 8'h25)? 32'h2cb59e09
	         : (byte_in == 8'h26)? 32'h1421b99b
	         : (byte_in == 8'h27)? 32'h2798798b
	         : (byte_in == 8'h28)? 32'h6508f6be
	         : (byte_in == 8'h29)? 32'h56b136ae
	         : (byte_in == 8'h2a)? 32'h6e25113c
	         : (byte_in == 8'h2b)? 32'h5d9cd12c
	         : (byte_in == 8'h2c)? 32'h3aef510d
	         : (byte_in == 8'h2d)? 32'h0956911d
	         : (byte_in == 8'h2e)? 32'h31c2b68f
	         : (byte_in == 8'h2f)? 32'h027b769f
	         : (byte_in == 8'h30)? 32'hcc9d76dd
	         : (byte_in == 8'h31)? 32'hff24b6cd
	         : (byte_in == 8'h32)? 32'hc7b0915f
	         : (byte_in == 8'h33)? 32'hf409514f
	         : (byte_in == 8'h34)? 32'h937ad16e
	         : (byte_in == 8'h35)? 32'ha0c3117e
	         : (byte_in == 8'h36)? 32'h985736ec
	         : (byte_in == 8'h37)? 32'habeef6fc
	         : (byte_in == 8'h38)? 32'he97e79c9
	         : (byte_in == 8'h39)? 32'hdac7b9d9
	         : (byte_in == 8'h3a)? 32'he2539e4b
	         : (byte_in == 8'h3b)? 32'hd1ea5e5b
	         : (byte_in == 8'h3c)? 32'hb699de7a
	         : (byte_in == 8'h3d)? 32'h85201e6a
	         : (byte_in == 8'h3e)? 32'hbdb439f8
	         : (byte_in == 8'h3f)? 32'h8e0df9e8
	         : (byte_in == 8'h40)? 32'h2079397d
	         : (byte_in == 8'h41)? 32'h13c0f96d
	         : (byte_in == 8'h42)? 32'h2b54deff
	         : (byte_in == 8'h43)? 32'h18ed1eef
	         : (byte_in == 8'h44)? 32'h7f9e9ece
	         : (byte_in == 8'h45)? 32'h4c275ede
	         : (byte_in == 8'h46)? 32'h74b3794c
	         : (byte_in == 8'h47)? 32'h470ab95c
	         : (byte_in == 8'h48)? 32'h059a3669
	         : (byte_in == 8'h49)? 32'h3623f679
	         : (byte_in == 8'h4a)? 32'h0eb7d1eb
	         : (byte_in == 8'h4b)? 32'h3d0e11fb
	         : (byte_in == 8'h4c)? 32'h5a7d91da
	         : (byte_in == 8'h4d)? 32'h69c451ca
	         : (byte_in == 8'h4e)? 32'h51507658
	         : (byte_in == 8'h4f)? 32'h62e9b648
	         : (byte_in == 8'h50)? 32'hac0fb60a
	         : (byte_in == 8'h51)? 32'h9fb6761a
	         : (byte_in == 8'h52)? 32'ha7225188
	         : (byte_in == 8'h53)? 32'h949b9198
	         : (byte_in == 8'h54)? 32'hf3e811b9
	         : (byte_in == 8'h55)? 32'hc051d1a9
	         : (byte_in == 8'h56)? 32'hf8c5f63b
	         : (byte_in == 8'h57)? 32'hcb7c362b
	         : (byte_in == 8'h58)? 32'h89ecb91e
	         : (byte_in == 8'h59)? 32'hba55790e
	         : (byte_in == 8'h5a)? 32'h82c15e9c
	         : (byte_in == 8'h5b)? 32'hb1789e8c
	         : (byte_in == 8'h5c)? 32'hd60b1ead
	         : (byte_in == 8'h5d)? 32'he5b2debd
	         : (byte_in == 8'h5e)? 32'hdd26f92f
	         : (byte_in == 8'h5f)? 32'hee9f393f
	         : (byte_in == 8'h60)? 32'h6092c0d7
	         : (byte_in == 8'h61)? 32'h532b00c7
	         : (byte_in == 8'h62)? 32'h6bbf2755
	         : (byte_in == 8'h63)? 32'h5806e745
	         : (byte_in == 8'h64)? 32'h3f756764
	         : (byte_in == 8'h65)? 32'h0ccca774
	         : (byte_in == 8'h66)? 32'h345880e6
	         : (byte_in == 8'h67)? 32'h07e140f6
	         : (byte_in == 8'h68)? 32'h4571cfc3
	         : (byte_in == 8'h69)? 32'h76c80fd3
	         : (byte_in == 8'h6a)? 32'h4e5c2841
	         : (byte_in == 8'h6b)? 32'h7de5e851
	         : (byte_in == 8'h6c)? 32'h1a966870
	         : (byte_in == 8'h6d)? 32'h292fa860
	         : (byte_in == 8'h6e)? 32'h11bb8ff2
	         : (byte_in == 8'h6f)? 32'h22024fe2
	         : (byte_in == 8'h70)? 32'hece44fa0
	         : (byte_in == 8'h71)? 32'hdf5d8fb0
	         : (byte_in == 8'h72)? 32'he7c9a822
	         : (byte_in == 8'h73)? 32'hd4706832
	         : (byte_in == 8'h74)? 32'hb303e813
	         : (byte_in == 8'h75)? 32'h80ba2803
	         : (byte_in == 8'h76)? 32'hb82e0f91
	         : (byte_in == 8'h77)? 32'h8b97cf81
	         : (byte_in == 8'h78)? 32'hc90740b4
	         : (byte_in == 8'h79)? 32'hfabe80a4
	         : (byte_in == 8'h7a)? 32'hc22aa736
	         : (byte_in == 8'h7b)? 32'hf1936726
	         : (byte_in == 8'h7c)? 32'h96e0e707
	         : (byte_in == 8'h7d)? 32'ha5592717
	         : (byte_in == 8'h7e)? 32'h9dcd0085
	         : (byte_in == 8'h7f)? 32'hae74c095
	         : (byte_in == 8'h80)? 32'hb26e3344
	         : (byte_in == 8'h81)? 32'h81d7f354
	         : (byte_in == 8'h82)? 32'hb943d4c6
	         : (byte_in == 8'h83)? 32'h8afa14d6
	         : (byte_in == 8'h84)? 32'hed8994f7
	         : (byte_in == 8'h85)? 32'hde3054e7
	         : (byte_in == 8'h86)? 32'he6a47375
	         : (byte_in == 8'h87)? 32'hd51db365
	         : (byte_in == 8'h88)? 32'h978d3c50
	         : (byte_in == 8'h89)? 32'ha434fc40
	         : (byte_in == 8'h8a)? 32'h9ca0dbd2
	         : (byte_in == 8'h8b)? 32'haf191bc2
	         : (byte_in == 8'h8c)? 32'hc86a9be3
	         : (byte_in == 8'h8d)? 32'hfbd35bf3
	         : (byte_in == 8'h8e)? 32'hc3477c61
	         : (byte_in == 8'h8f)? 32'hf0febc71
	         : (byte_in == 8'h90)? 32'h3e18bc33
	         : (byte_in == 8'h91)? 32'h0da17c23
	         : (byte_in == 8'h92)? 32'h35355bb1
	         : (byte_in == 8'h93)? 32'h068c9ba1
	         : (byte_in == 8'h94)? 32'h61ff1b80
	         : (byte_in == 8'h95)? 32'h5246db90
	         : (byte_in == 8'h96)? 32'h6ad2fc02
	         : (byte_in == 8'h97)? 32'h596b3c12
	         : (byte_in == 8'h98)? 32'h1bfbb327
	         : (byte_in == 8'h99)? 32'h28427337
	         : (byte_in == 8'h9a)? 32'h10d654a5
	         : (byte_in == 8'h9b)? 32'h236f94b5
	         : (byte_in == 8'h9c)? 32'h441c1494
	         : (byte_in == 8'h9d)? 32'h77a5d484
	         : (byte_in == 8'h9e)? 32'h4f31f316
	         : (byte_in == 8'h9f)? 32'h7c883306
	         : (byte_in == 8'ha0)? 32'hf285caee
	         : (byte_in == 8'ha1)? 32'hc13c0afe
	         : (byte_in == 8'ha2)? 32'hf9a82d6c
	         : (byte_in == 8'ha3)? 32'hca11ed7c
	         : (byte_in == 8'ha4)? 32'had626d5d
	         : (byte_in == 8'ha5)? 32'h9edbad4d
	         : (byte_in == 8'ha6)? 32'ha64f8adf
	         : (byte_in == 8'ha7)? 32'h95f64acf
	         : (byte_in == 8'ha8)? 32'hd766c5fa
	         : (byte_in == 8'ha9)? 32'he4df05ea
	         : (byte_in == 8'haa)? 32'hdc4b2278
	         : (byte_in == 8'hab)? 32'heff2e268
	         : (byte_in == 8'hac)? 32'h88816249
	         : (byte_in == 8'had)? 32'hbb38a259
	         : (byte_in == 8'hae)? 32'h83ac85cb
	         : (byte_in == 8'haf)? 32'hb01545db
	         : (byte_in == 8'hb0)? 32'h7ef34599
	         : (byte_in == 8'hb1)? 32'h4d4a8589
	         : (byte_in == 8'hb2)? 32'h75dea21b
	         : (byte_in == 8'hb3)? 32'h4667620b
	         : (byte_in == 8'hb4)? 32'h2114e22a
	         : (byte_in == 8'hb5)? 32'h12ad223a
	         : (byte_in == 8'hb6)? 32'h2a3905a8
	         : (byte_in == 8'hb7)? 32'h1980c5b8
	         : (byte_in == 8'hb8)? 32'h5b104a8d
	         : (byte_in == 8'hb9)? 32'h68a98a9d
	         : (byte_in == 8'hba)? 32'h503dad0f
	         : (byte_in == 8'hbb)? 32'h63846d1f
	         : (byte_in == 8'hbc)? 32'h04f7ed3e
	         : (byte_in == 8'hbd)? 32'h374e2d2e
	         : (byte_in == 8'hbe)? 32'h0fda0abc
	         : (byte_in == 8'hbf)? 32'h3c63caac
	         : (byte_in == 8'hc0)? 32'h92170a39
	         : (byte_in == 8'hc1)? 32'ha1aeca29
	         : (byte_in == 8'hc2)? 32'h993aedbb
	         : (byte_in == 8'hc3)? 32'haa832dab
	         : (byte_in == 8'hc4)? 32'hcdf0ad8a
	         : (byte_in == 8'hc5)? 32'hfe496d9a
	         : (byte_in == 8'hc6)? 32'hc6dd4a08
	         : (byte_in == 8'hc7)? 32'hf5648a18
	         : (byte_in == 8'hc8)? 32'hb7f4052d
	         : (byte_in == 8'hc9)? 32'h844dc53d
	         : (byte_in == 8'hca)? 32'hbcd9e2af
	         : (byte_in == 8'hcb)? 32'h8f6022bf
	         : (byte_in == 8'hcc)? 32'he813a29e
	         : (byte_in == 8'hcd)? 32'hdbaa628e
	         : (byte_in == 8'hce)? 32'he33e451c
	         : (byte_in == 8'hcf)? 32'hd087850c
	         : (byte_in == 8'hd0)? 32'h1e61854e
	         : (byte_in == 8'hd1)? 32'h2dd8455e
	         : (byte_in == 8'hd2)? 32'h154c62cc
	         : (byte_in == 8'hd3)? 32'h26f5a2dc
	         : (byte_in == 8'hd4)? 32'h418622fd
	         : (byte_in == 8'hd5)? 32'h723fe2ed
	         : (byte_in == 8'hd6)? 32'h4aabc57f
	         : (byte_in == 8'hd7)? 32'h7912056f
	         : (byte_in == 8'hd8)? 32'h3b828a5a
	         : (byte_in == 8'hd9)? 32'h083b4a4a
	         : (byte_in == 8'hda)? 32'h30af6dd8
	         : (byte_in == 8'hdb)? 32'h0316adc8
	         : (byte_in == 8'hdc)? 32'h64652de9
	         : (byte_in == 8'hdd)? 32'h57dcedf9
	         : (byte_in == 8'hde)? 32'h6f48ca6b
	         : (byte_in == 8'hdf)? 32'h5cf10a7b
	         : (byte_in == 8'he0)? 32'hd2fcf393
	         : (byte_in == 8'he1)? 32'he1453383
	         : (byte_in == 8'he2)? 32'hd9d11411
	         : (byte_in == 8'he3)? 32'hea68d401
	         : (byte_in == 8'he4)? 32'h8d1b5420
	         : (byte_in == 8'he5)? 32'hbea29430
	         : (byte_in == 8'he6)? 32'h8636b3a2
	         : (byte_in == 8'he7)? 32'hb58f73b2
	         : (byte_in == 8'he8)? 32'hf71ffc87
	         : (byte_in == 8'he9)? 32'hc4a63c97
	         : (byte_in == 8'hea)? 32'hfc321b05
	         : (byte_in == 8'heb)? 32'hcf8bdb15
	         : (byte_in == 8'hec)? 32'ha8f85b34
	         : (byte_in == 8'hed)? 32'h9b419b24
	         : (byte_in == 8'hee)? 32'ha3d5bcb6
	         : (byte_in == 8'hef)? 32'h906c7ca6
	         : (byte_in == 8'hf0)? 32'h5e8a7ce4
	         : (byte_in == 8'hf1)? 32'h6d33bcf4
	         : (byte_in == 8'hf2)? 32'h55a79b66
	         : (byte_in == 8'hf3)? 32'h661e5b76
	         : (byte_in == 8'hf4)? 32'h016ddb57
	         : (byte_in == 8'hf5)? 32'h32d41b47
	         : (byte_in == 8'hf6)? 32'h0a403cd5
	         : (byte_in == 8'hf7)? 32'h39f9fcc5
	         : (byte_in == 8'hf8)? 32'h7b6973f0
	         : (byte_in == 8'hf9)? 32'h48d0b3e0
	         : (byte_in == 8'hfa)? 32'h70449472
	         : (byte_in == 8'hfb)? 32'h43fd5462
	         : (byte_in == 8'hfc)? 32'h248ed443
	         : (byte_in == 8'hfd)? 32'h17371453
	         : (byte_in == 8'hfe)? 32'h2fa333c1
	         :                     32'h1c1af3d1;

endmodule
//}}}

module TABLE5(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h40f372fb
	         : (byte_in == 8'h02)? 32'h64dd6689
	         : (byte_in == 8'h03)? 32'h242e1472
	         : (byte_in == 8'h04)? 32'h81e7e5f6
	         : (byte_in == 8'h05)? 32'hc114970d
	         : (byte_in == 8'h06)? 32'he53a837f
	         : (byte_in == 8'h07)? 32'ha5c9f184
	         : (byte_in == 8'h08)? 32'hc9bacd12
	         : (byte_in == 8'h09)? 32'h8949bfe9
	         : (byte_in == 8'h0a)? 32'had67ab9b
	         : (byte_in == 8'h0b)? 32'hed94d960
	         : (byte_in == 8'h0c)? 32'h485d28e4
	         : (byte_in == 8'h0d)? 32'h08ae5a1f
	         : (byte_in == 8'h0e)? 32'h2c804e6d
	         : (byte_in == 8'h0f)? 32'h6c733c96
	         : (byte_in == 8'h10)? 32'h3b5bec7e
	         : (byte_in == 8'h11)? 32'h7ba89e85
	         : (byte_in == 8'h12)? 32'h5f868af7
	         : (byte_in == 8'h13)? 32'h1f75f80c
	         : (byte_in == 8'h14)? 32'hbabc0988
	         : (byte_in == 8'h15)? 32'hfa4f7b73
	         : (byte_in == 8'h16)? 32'hde616f01
	         : (byte_in == 8'h17)? 32'h9e921dfa
	         : (byte_in == 8'h18)? 32'hf2e1216c
	         : (byte_in == 8'h19)? 32'hb2125397
	         : (byte_in == 8'h1a)? 32'h963c47e5
	         : (byte_in == 8'h1b)? 32'hd6cf351e
	         : (byte_in == 8'h1c)? 32'h7306c49a
	         : (byte_in == 8'h1d)? 32'h33f5b661
	         : (byte_in == 8'h1e)? 32'h17dba213
	         : (byte_in == 8'h1f)? 32'h5728d0e8
	         : (byte_in == 8'h20)? 32'ha0cd5a34
	         : (byte_in == 8'h21)? 32'he03e28cf
	         : (byte_in == 8'h22)? 32'hc4103cbd
	         : (byte_in == 8'h23)? 32'h84e34e46
	         : (byte_in == 8'h24)? 32'h212abfc2
	         : (byte_in == 8'h25)? 32'h61d9cd39
	         : (byte_in == 8'h26)? 32'h45f7d94b
	         : (byte_in == 8'h27)? 32'h0504abb0
	         : (byte_in == 8'h28)? 32'h69779726
	         : (byte_in == 8'h29)? 32'h2984e5dd
	         : (byte_in == 8'h2a)? 32'h0daaf1af
	         : (byte_in == 8'h2b)? 32'h4d598354
	         : (byte_in == 8'h2c)? 32'he89072d0
	         : (byte_in == 8'h2d)? 32'ha863002b
	         : (byte_in == 8'h2e)? 32'h8c4d1459
	         : (byte_in == 8'h2f)? 32'hccbe66a2
	         : (byte_in == 8'h30)? 32'h9b96b64a
	         : (byte_in == 8'h31)? 32'hdb65c4b1
	         : (byte_in == 8'h32)? 32'hff4bd0c3
	         : (byte_in == 8'h33)? 32'hbfb8a238
	         : (byte_in == 8'h34)? 32'h1a7153bc
	         : (byte_in == 8'h35)? 32'h5a822147
	         : (byte_in == 8'h36)? 32'h7eac3535
	         : (byte_in == 8'h37)? 32'h3e5f47ce
	         : (byte_in == 8'h38)? 32'h522c7b58
	         : (byte_in == 8'h39)? 32'h12df09a3
	         : (byte_in == 8'h3a)? 32'h36f11dd1
	         : (byte_in == 8'h3b)? 32'h76026f2a
	         : (byte_in == 8'h3c)? 32'hd3cb9eae
	         : (byte_in == 8'h3d)? 32'h9338ec55
	         : (byte_in == 8'h3e)? 32'hb716f827
	         : (byte_in == 8'h3f)? 32'hf7e58adc
	         : (byte_in == 8'h40)? 32'h450f18ec
	         : (byte_in == 8'h41)? 32'h05fc6a17
	         : (byte_in == 8'h42)? 32'h21d27e65
	         : (byte_in == 8'h43)? 32'h61210c9e
	         : (byte_in == 8'h44)? 32'hc4e8fd1a
	         : (byte_in == 8'h45)? 32'h841b8fe1
	         : (byte_in == 8'h46)? 32'ha0359b93
	         : (byte_in == 8'h47)? 32'he0c6e968
	         : (byte_in == 8'h48)? 32'h8cb5d5fe
	         : (byte_in == 8'h49)? 32'hcc46a705
	         : (byte_in == 8'h4a)? 32'he868b377
	         : (byte_in == 8'h4b)? 32'ha89bc18c
	         : (byte_in == 8'h4c)? 32'h0d523008
	         : (byte_in == 8'h4d)? 32'h4da142f3
	         : (byte_in == 8'h4e)? 32'h698f5681
	         : (byte_in == 8'h4f)? 32'h297c247a
	         : (byte_in == 8'h50)? 32'h7e54f492
	         : (byte_in == 8'h51)? 32'h3ea78669
	         : (byte_in == 8'h52)? 32'h1a89921b
	         : (byte_in == 8'h53)? 32'h5a7ae0e0
	         : (byte_in == 8'h54)? 32'hffb31164
	         : (byte_in == 8'h55)? 32'hbf40639f
	         : (byte_in == 8'h56)? 32'h9b6e77ed
	         : (byte_in == 8'h57)? 32'hdb9d0516
	         : (byte_in == 8'h58)? 32'hb7ee3980
	         : (byte_in == 8'h59)? 32'hf71d4b7b
	         : (byte_in == 8'h5a)? 32'hd3335f09
	         : (byte_in == 8'h5b)? 32'h93c02df2
	         : (byte_in == 8'h5c)? 32'h3609dc76
	         : (byte_in == 8'h5d)? 32'h76faae8d
	         : (byte_in == 8'h5e)? 32'h52d4baff
	         : (byte_in == 8'h5f)? 32'h1227c804
	         : (byte_in == 8'h60)? 32'he5c242d8
	         : (byte_in == 8'h61)? 32'ha5313023
	         : (byte_in == 8'h62)? 32'h811f2451
	         : (byte_in == 8'h63)? 32'hc1ec56aa
	         : (byte_in == 8'h64)? 32'h6425a72e
	         : (byte_in == 8'h65)? 32'h24d6d5d5
	         : (byte_in == 8'h66)? 32'h00f8c1a7
	         : (byte_in == 8'h67)? 32'h400bb35c
	         : (byte_in == 8'h68)? 32'h2c788fca
	         : (byte_in == 8'h69)? 32'h6c8bfd31
	         : (byte_in == 8'h6a)? 32'h48a5e943
	         : (byte_in == 8'h6b)? 32'h08569bb8
	         : (byte_in == 8'h6c)? 32'had9f6a3c
	         : (byte_in == 8'h6d)? 32'hed6c18c7
	         : (byte_in == 8'h6e)? 32'hc9420cb5
	         : (byte_in == 8'h6f)? 32'h89b17e4e
	         : (byte_in == 8'h70)? 32'hde99aea6
	         : (byte_in == 8'h71)? 32'h9e6adc5d
	         : (byte_in == 8'h72)? 32'hba44c82f
	         : (byte_in == 8'h73)? 32'hfab7bad4
	         : (byte_in == 8'h74)? 32'h5f7e4b50
	         : (byte_in == 8'h75)? 32'h1f8d39ab
	         : (byte_in == 8'h76)? 32'h3ba32dd9
	         : (byte_in == 8'h77)? 32'h7b505f22
	         : (byte_in == 8'h78)? 32'h172363b4
	         : (byte_in == 8'h79)? 32'h57d0114f
	         : (byte_in == 8'h7a)? 32'h73fe053d
	         : (byte_in == 8'h7b)? 32'h330d77c6
	         : (byte_in == 8'h7c)? 32'h96c48642
	         : (byte_in == 8'h7d)? 32'hd637f4b9
	         : (byte_in == 8'h7e)? 32'hf219e0cb
	         : (byte_in == 8'h7f)? 32'hb2ea9230
	         : (byte_in == 8'h80)? 32'h4ab753eb
	         : (byte_in == 8'h81)? 32'h0a442110
	         : (byte_in == 8'h82)? 32'h2e6a3562
	         : (byte_in == 8'h83)? 32'h6e994799
	         : (byte_in == 8'h84)? 32'hcb50b61d
	         : (byte_in == 8'h85)? 32'h8ba3c4e6
	         : (byte_in == 8'h86)? 32'haf8dd094
	         : (byte_in == 8'h87)? 32'hef7ea26f
	         : (byte_in == 8'h88)? 32'h830d9ef9
	         : (byte_in == 8'h89)? 32'hc3feec02
	         : (byte_in == 8'h8a)? 32'he7d0f870
	         : (byte_in == 8'h8b)? 32'ha7238a8b
	         : (byte_in == 8'h8c)? 32'h02ea7b0f
	         : (byte_in == 8'h8d)? 32'h421909f4
	         : (byte_in == 8'h8e)? 32'h66371d86
	         : (byte_in == 8'h8f)? 32'h26c46f7d
	         : (byte_in == 8'h90)? 32'h71ecbf95
	         : (byte_in == 8'h91)? 32'h311fcd6e
	         : (byte_in == 8'h92)? 32'h1531d91c
	         : (byte_in == 8'h93)? 32'h55c2abe7
	         : (byte_in == 8'h94)? 32'hf00b5a63
	         : (byte_in == 8'h95)? 32'hb0f82898
	         : (byte_in == 8'h96)? 32'h94d63cea
	         : (byte_in == 8'h97)? 32'hd4254e11
	         : (byte_in == 8'h98)? 32'hb8567287
	         : (byte_in == 8'h99)? 32'hf8a5007c
	         : (byte_in == 8'h9a)? 32'hdc8b140e
	         : (byte_in == 8'h9b)? 32'h9c7866f5
	         : (byte_in == 8'h9c)? 32'h39b19771
	         : (byte_in == 8'h9d)? 32'h7942e58a
	         : (byte_in == 8'h9e)? 32'h5d6cf1f8
	         : (byte_in == 8'h9f)? 32'h1d9f8303
	         : (byte_in == 8'ha0)? 32'hea7a09df
	         : (byte_in == 8'ha1)? 32'haa897b24
	         : (byte_in == 8'ha2)? 32'h8ea76f56
	         : (byte_in == 8'ha3)? 32'hce541dad
	         : (byte_in == 8'ha4)? 32'h6b9dec29
	         : (byte_in == 8'ha5)? 32'h2b6e9ed2
	         : (byte_in == 8'ha6)? 32'h0f408aa0
	         : (byte_in == 8'ha7)? 32'h4fb3f85b
	         : (byte_in == 8'ha8)? 32'h23c0c4cd
	         : (byte_in == 8'ha9)? 32'h6333b636
	         : (byte_in == 8'haa)? 32'h471da244
	         : (byte_in == 8'hab)? 32'h07eed0bf
	         : (byte_in == 8'hac)? 32'ha227213b
	         : (byte_in == 8'had)? 32'he2d453c0
	         : (byte_in == 8'hae)? 32'hc6fa47b2
	         : (byte_in == 8'haf)? 32'h86093549
	         : (byte_in == 8'hb0)? 32'hd121e5a1
	         : (byte_in == 8'hb1)? 32'h91d2975a
	         : (byte_in == 8'hb2)? 32'hb5fc8328
	         : (byte_in == 8'hb3)? 32'hf50ff1d3
	         : (byte_in == 8'hb4)? 32'h50c60057
	         : (byte_in == 8'hb5)? 32'h103572ac
	         : (byte_in == 8'hb6)? 32'h341b66de
	         : (byte_in == 8'hb7)? 32'h74e81425
	         : (byte_in == 8'hb8)? 32'h189b28b3
	         : (byte_in == 8'hb9)? 32'h58685a48
	         : (byte_in == 8'hba)? 32'h7c464e3a
	         : (byte_in == 8'hbb)? 32'h3cb53cc1
	         : (byte_in == 8'hbc)? 32'h997ccd45
	         : (byte_in == 8'hbd)? 32'hd98fbfbe
	         : (byte_in == 8'hbe)? 32'hfda1abcc
	         : (byte_in == 8'hbf)? 32'hbd52d937
	         : (byte_in == 8'hc0)? 32'h0fb84b07
	         : (byte_in == 8'hc1)? 32'h4f4b39fc
	         : (byte_in == 8'hc2)? 32'h6b652d8e
	         : (byte_in == 8'hc3)? 32'h2b965f75
	         : (byte_in == 8'hc4)? 32'h8e5faef1
	         : (byte_in == 8'hc5)? 32'hceacdc0a
	         : (byte_in == 8'hc6)? 32'hea82c878
	         : (byte_in == 8'hc7)? 32'haa71ba83
	         : (byte_in == 8'hc8)? 32'hc6028615
	         : (byte_in == 8'hc9)? 32'h86f1f4ee
	         : (byte_in == 8'hca)? 32'ha2dfe09c
	         : (byte_in == 8'hcb)? 32'he22c9267
	         : (byte_in == 8'hcc)? 32'h47e563e3
	         : (byte_in == 8'hcd)? 32'h07161118
	         : (byte_in == 8'hce)? 32'h2338056a
	         : (byte_in == 8'hcf)? 32'h63cb7791
	         : (byte_in == 8'hd0)? 32'h34e3a779
	         : (byte_in == 8'hd1)? 32'h7410d582
	         : (byte_in == 8'hd2)? 32'h503ec1f0
	         : (byte_in == 8'hd3)? 32'h10cdb30b
	         : (byte_in == 8'hd4)? 32'hb504428f
	         : (byte_in == 8'hd5)? 32'hf5f73074
	         : (byte_in == 8'hd6)? 32'hd1d92406
	         : (byte_in == 8'hd7)? 32'h912a56fd
	         : (byte_in == 8'hd8)? 32'hfd596a6b
	         : (byte_in == 8'hd9)? 32'hbdaa1890
	         : (byte_in == 8'hda)? 32'h99840ce2
	         : (byte_in == 8'hdb)? 32'hd9777e19
	         : (byte_in == 8'hdc)? 32'h7cbe8f9d
	         : (byte_in == 8'hdd)? 32'h3c4dfd66
	         : (byte_in == 8'hde)? 32'h1863e914
	         : (byte_in == 8'hdf)? 32'h58909bef
	         : (byte_in == 8'he0)? 32'haf751133
	         : (byte_in == 8'he1)? 32'hef8663c8
	         : (byte_in == 8'he2)? 32'hcba877ba
	         : (byte_in == 8'he3)? 32'h8b5b0541
	         : (byte_in == 8'he4)? 32'h2e92f4c5
	         : (byte_in == 8'he5)? 32'h6e61863e
	         : (byte_in == 8'he6)? 32'h4a4f924c
	         : (byte_in == 8'he7)? 32'h0abce0b7
	         : (byte_in == 8'he8)? 32'h66cfdc21
	         : (byte_in == 8'he9)? 32'h263caeda
	         : (byte_in == 8'hea)? 32'h0212baa8
	         : (byte_in == 8'heb)? 32'h42e1c853
	         : (byte_in == 8'hec)? 32'he72839d7
	         : (byte_in == 8'hed)? 32'ha7db4b2c
	         : (byte_in == 8'hee)? 32'h83f55f5e
	         : (byte_in == 8'hef)? 32'hc3062da5
	         : (byte_in == 8'hf0)? 32'h942efd4d
	         : (byte_in == 8'hf1)? 32'hd4dd8fb6
	         : (byte_in == 8'hf2)? 32'hf0f39bc4
	         : (byte_in == 8'hf3)? 32'hb000e93f
	         : (byte_in == 8'hf4)? 32'h15c918bb
	         : (byte_in == 8'hf5)? 32'h553a6a40
	         : (byte_in == 8'hf6)? 32'h71147e32
	         : (byte_in == 8'hf7)? 32'h31e70cc9
	         : (byte_in == 8'hf8)? 32'h5d94305f
	         : (byte_in == 8'hf9)? 32'h1d6742a4
	         : (byte_in == 8'hfa)? 32'h394956d6
	         : (byte_in == 8'hfb)? 32'h79ba242d
	         : (byte_in == 8'hfc)? 32'hdc73d5a9
	         : (byte_in == 8'hfd)? 32'h9c80a752
	         : (byte_in == 8'hfe)? 32'hb8aeb320
	         :                     32'hf85dc1db;

endmodule
//}}}

module TABLE6(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h8a1f31d8
	         : (byte_in == 8'h02)? 32'h956fa7d6
	         : (byte_in == 8'h03)? 32'h1f70960e
	         : (byte_in == 8'h04)? 32'h1f128433
	         : (byte_in == 8'h05)? 32'h950db5eb
	         : (byte_in == 8'h06)? 32'h8a7d23e5
	         : (byte_in == 8'h07)? 32'h0062123d
	         : (byte_in == 8'h08)? 32'h124b683e
	         : (byte_in == 8'h09)? 32'h985459e6
	         : (byte_in == 8'h0a)? 32'h8724cfe8
	         : (byte_in == 8'h0b)? 32'h0d3bfe30
	         : (byte_in == 8'h0c)? 32'h0d59ec0d
	         : (byte_in == 8'h0d)? 32'h8746ddd5
	         : (byte_in == 8'h0e)? 32'h98364bdb
	         : (byte_in == 8'h0f)? 32'h12297a03
	         : (byte_in == 8'h10)? 32'h0d9dc877
	         : (byte_in == 8'h11)? 32'h8782f9af
	         : (byte_in == 8'h12)? 32'h98f26fa1
	         : (byte_in == 8'h13)? 32'h12ed5e79
	         : (byte_in == 8'h14)? 32'h128f4c44
	         : (byte_in == 8'h15)? 32'h98907d9c
	         : (byte_in == 8'h16)? 32'h87e0eb92
	         : (byte_in == 8'h17)? 32'h0dffda4a
	         : (byte_in == 8'h18)? 32'h1fd6a049
	         : (byte_in == 8'h19)? 32'h95c99191
	         : (byte_in == 8'h1a)? 32'h8ab9079f
	         : (byte_in == 8'h1b)? 32'h00a63647
	         : (byte_in == 8'h1c)? 32'h00c4247a
	         : (byte_in == 8'h1d)? 32'h8adb15a2
	         : (byte_in == 8'h1e)? 32'h95ab83ac
	         : (byte_in == 8'h1f)? 32'h1fb4b274
	         : (byte_in == 8'h20)? 32'h2fba37ff
	         : (byte_in == 8'h21)? 32'ha5a50627
	         : (byte_in == 8'h22)? 32'hbad59029
	         : (byte_in == 8'h23)? 32'h30caa1f1
	         : (byte_in == 8'h24)? 32'h30a8b3cc
	         : (byte_in == 8'h25)? 32'hbab78214
	         : (byte_in == 8'h26)? 32'ha5c7141a
	         : (byte_in == 8'h27)? 32'h2fd825c2
	         : (byte_in == 8'h28)? 32'h3df15fc1
	         : (byte_in == 8'h29)? 32'hb7ee6e19
	         : (byte_in == 8'h2a)? 32'ha89ef817
	         : (byte_in == 8'h2b)? 32'h2281c9cf
	         : (byte_in == 8'h2c)? 32'h22e3dbf2
	         : (byte_in == 8'h2d)? 32'ha8fcea2a
	         : (byte_in == 8'h2e)? 32'hb78c7c24
	         : (byte_in == 8'h2f)? 32'h3d934dfc
	         : (byte_in == 8'h30)? 32'h2227ff88
	         : (byte_in == 8'h31)? 32'ha838ce50
	         : (byte_in == 8'h32)? 32'hb748585e
	         : (byte_in == 8'h33)? 32'h3d576986
	         : (byte_in == 8'h34)? 32'h3d357bbb
	         : (byte_in == 8'h35)? 32'hb72a4a63
	         : (byte_in == 8'h36)? 32'ha85adc6d
	         : (byte_in == 8'h37)? 32'h2245edb5
	         : (byte_in == 8'h38)? 32'h306c97b6
	         : (byte_in == 8'h39)? 32'hba73a66e
	         : (byte_in == 8'h3a)? 32'ha5033060
	         : (byte_in == 8'h3b)? 32'h2f1c01b8
	         : (byte_in == 8'h3c)? 32'h2f7e1385
	         : (byte_in == 8'h3d)? 32'ha561225d
	         : (byte_in == 8'h3e)? 32'hba11b453
	         : (byte_in == 8'h3f)? 32'h300e858b
	         : (byte_in == 8'h40)? 32'h288350fe
	         : (byte_in == 8'h41)? 32'ha29c6126
	         : (byte_in == 8'h42)? 32'hbdecf728
	         : (byte_in == 8'h43)? 32'h37f3c6f0
	         : (byte_in == 8'h44)? 32'h3791d4cd
	         : (byte_in == 8'h45)? 32'hbd8ee515
	         : (byte_in == 8'h46)? 32'ha2fe731b
	         : (byte_in == 8'h47)? 32'h28e142c3
	         : (byte_in == 8'h48)? 32'h3ac838c0
	         : (byte_in == 8'h49)? 32'hb0d70918
	         : (byte_in == 8'h4a)? 32'hafa79f16
	         : (byte_in == 8'h4b)? 32'h25b8aece
	         : (byte_in == 8'h4c)? 32'h25dabcf3
	         : (byte_in == 8'h4d)? 32'hafc58d2b
	         : (byte_in == 8'h4e)? 32'hb0b51b25
	         : (byte_in == 8'h4f)? 32'h3aaa2afd
	         : (byte_in == 8'h50)? 32'h251e9889
	         : (byte_in == 8'h51)? 32'haf01a951
	         : (byte_in == 8'h52)? 32'hb0713f5f
	         : (byte_in == 8'h53)? 32'h3a6e0e87
	         : (byte_in == 8'h54)? 32'h3a0c1cba
	         : (byte_in == 8'h55)? 32'hb0132d62
	         : (byte_in == 8'h56)? 32'haf63bb6c
	         : (byte_in == 8'h57)? 32'h257c8ab4
	         : (byte_in == 8'h58)? 32'h3755f0b7
	         : (byte_in == 8'h59)? 32'hbd4ac16f
	         : (byte_in == 8'h5a)? 32'ha23a5761
	         : (byte_in == 8'h5b)? 32'h282566b9
	         : (byte_in == 8'h5c)? 32'h28477484
	         : (byte_in == 8'h5d)? 32'ha258455c
	         : (byte_in == 8'h5e)? 32'hbd28d352
	         : (byte_in == 8'h5f)? 32'h3737e28a
	         : (byte_in == 8'h60)? 32'h07396701
	         : (byte_in == 8'h61)? 32'h8d2656d9
	         : (byte_in == 8'h62)? 32'h9256c0d7
	         : (byte_in == 8'h63)? 32'h1849f10f
	         : (byte_in == 8'h64)? 32'h182be332
	         : (byte_in == 8'h65)? 32'h9234d2ea
	         : (byte_in == 8'h66)? 32'h8d4444e4
	         : (byte_in == 8'h67)? 32'h075b753c
	         : (byte_in == 8'h68)? 32'h15720f3f
	         : (byte_in == 8'h69)? 32'h9f6d3ee7
	         : (byte_in == 8'h6a)? 32'h801da8e9
	         : (byte_in == 8'h6b)? 32'h0a029931
	         : (byte_in == 8'h6c)? 32'h0a608b0c
	         : (byte_in == 8'h6d)? 32'h807fbad4
	         : (byte_in == 8'h6e)? 32'h9f0f2cda
	         : (byte_in == 8'h6f)? 32'h15101d02
	         : (byte_in == 8'h70)? 32'h0aa4af76
	         : (byte_in == 8'h71)? 32'h80bb9eae
	         : (byte_in == 8'h72)? 32'h9fcb08a0
	         : (byte_in == 8'h73)? 32'h15d43978
	         : (byte_in == 8'h74)? 32'h15b62b45
	         : (byte_in == 8'h75)? 32'h9fa91a9d
	         : (byte_in == 8'h76)? 32'h80d98c93
	         : (byte_in == 8'h77)? 32'h0ac6bd4b
	         : (byte_in == 8'h78)? 32'h18efc748
	         : (byte_in == 8'h79)? 32'h92f0f690
	         : (byte_in == 8'h7a)? 32'h8d80609e
	         : (byte_in == 8'h7b)? 32'h079f5146
	         : (byte_in == 8'h7c)? 32'h07fd437b
	         : (byte_in == 8'h7d)? 32'h8de272a3
	         : (byte_in == 8'h7e)? 32'h9292e4ad
	         : (byte_in == 8'h7f)? 32'h188dd575
	         : (byte_in == 8'h80)? 32'h5459887d
	         : (byte_in == 8'h81)? 32'hde46b9a5
	         : (byte_in == 8'h82)? 32'hc1362fab
	         : (byte_in == 8'h83)? 32'h4b291e73
	         : (byte_in == 8'h84)? 32'h4b4b0c4e
	         : (byte_in == 8'h85)? 32'hc1543d96
	         : (byte_in == 8'h86)? 32'hde24ab98
	         : (byte_in == 8'h87)? 32'h543b9a40
	         : (byte_in == 8'h88)? 32'h4612e043
	         : (byte_in == 8'h89)? 32'hcc0dd19b
	         : (byte_in == 8'h8a)? 32'hd37d4795
	         : (byte_in == 8'h8b)? 32'h5962764d
	         : (byte_in == 8'h8c)? 32'h59006470
	         : (byte_in == 8'h8d)? 32'hd31f55a8
	         : (byte_in == 8'h8e)? 32'hcc6fc3a6
	         : (byte_in == 8'h8f)? 32'h4670f27e
	         : (byte_in == 8'h90)? 32'h59c4400a
	         : (byte_in == 8'h91)? 32'hd3db71d2
	         : (byte_in == 8'h92)? 32'hccabe7dc
	         : (byte_in == 8'h93)? 32'h46b4d604
	         : (byte_in == 8'h94)? 32'h46d6c439
	         : (byte_in == 8'h95)? 32'hccc9f5e1
	         : (byte_in == 8'h96)? 32'hd3b963ef
	         : (byte_in == 8'h97)? 32'h59a65237
	         : (byte_in == 8'h98)? 32'h4b8f2834
	         : (byte_in == 8'h99)? 32'hc19019ec
	         : (byte_in == 8'h9a)? 32'hdee08fe2
	         : (byte_in == 8'h9b)? 32'h54ffbe3a
	         : (byte_in == 8'h9c)? 32'h549dac07
	         : (byte_in == 8'h9d)? 32'hde829ddf
	         : (byte_in == 8'h9e)? 32'hc1f20bd1
	         : (byte_in == 8'h9f)? 32'h4bed3a09
	         : (byte_in == 8'ha0)? 32'h7be3bf82
	         : (byte_in == 8'ha1)? 32'hf1fc8e5a
	         : (byte_in == 8'ha2)? 32'hee8c1854
	         : (byte_in == 8'ha3)? 32'h6493298c
	         : (byte_in == 8'ha4)? 32'h64f13bb1
	         : (byte_in == 8'ha5)? 32'heeee0a69
	         : (byte_in == 8'ha6)? 32'hf19e9c67
	         : (byte_in == 8'ha7)? 32'h7b81adbf
	         : (byte_in == 8'ha8)? 32'h69a8d7bc
	         : (byte_in == 8'ha9)? 32'he3b7e664
	         : (byte_in == 8'haa)? 32'hfcc7706a
	         : (byte_in == 8'hab)? 32'h76d841b2
	         : (byte_in == 8'hac)? 32'h76ba538f
	         : (byte_in == 8'had)? 32'hfca56257
	         : (byte_in == 8'hae)? 32'he3d5f459
	         : (byte_in == 8'haf)? 32'h69cac581
	         : (byte_in == 8'hb0)? 32'h767e77f5
	         : (byte_in == 8'hb1)? 32'hfc61462d
	         : (byte_in == 8'hb2)? 32'he311d023
	         : (byte_in == 8'hb3)? 32'h690ee1fb
	         : (byte_in == 8'hb4)? 32'h696cf3c6
	         : (byte_in == 8'hb5)? 32'he373c21e
	         : (byte_in == 8'hb6)? 32'hfc035410
	         : (byte_in == 8'hb7)? 32'h761c65c8
	         : (byte_in == 8'hb8)? 32'h64351fcb
	         : (byte_in == 8'hb9)? 32'hee2a2e13
	         : (byte_in == 8'hba)? 32'hf15ab81d
	         : (byte_in == 8'hbb)? 32'h7b4589c5
	         : (byte_in == 8'hbc)? 32'h7b279bf8
	         : (byte_in == 8'hbd)? 32'hf138aa20
	         : (byte_in == 8'hbe)? 32'hee483c2e
	         : (byte_in == 8'hbf)? 32'h64570df6
	         : (byte_in == 8'hc0)? 32'h7cdad883
	         : (byte_in == 8'hc1)? 32'hf6c5e95b
	         : (byte_in == 8'hc2)? 32'he9b57f55
	         : (byte_in == 8'hc3)? 32'h63aa4e8d
	         : (byte_in == 8'hc4)? 32'h63c85cb0
	         : (byte_in == 8'hc5)? 32'he9d76d68
	         : (byte_in == 8'hc6)? 32'hf6a7fb66
	         : (byte_in == 8'hc7)? 32'h7cb8cabe
	         : (byte_in == 8'hc8)? 32'h6e91b0bd
	         : (byte_in == 8'hc9)? 32'he48e8165
	         : (byte_in == 8'hca)? 32'hfbfe176b
	         : (byte_in == 8'hcb)? 32'h71e126b3
	         : (byte_in == 8'hcc)? 32'h7183348e
	         : (byte_in == 8'hcd)? 32'hfb9c0556
	         : (byte_in == 8'hce)? 32'he4ec9358
	         : (byte_in == 8'hcf)? 32'h6ef3a280
	         : (byte_in == 8'hd0)? 32'h714710f4
	         : (byte_in == 8'hd1)? 32'hfb58212c
	         : (byte_in == 8'hd2)? 32'he428b722
	         : (byte_in == 8'hd3)? 32'h6e3786fa
	         : (byte_in == 8'hd4)? 32'h6e5594c7
	         : (byte_in == 8'hd5)? 32'he44aa51f
	         : (byte_in == 8'hd6)? 32'hfb3a3311
	         : (byte_in == 8'hd7)? 32'h712502c9
	         : (byte_in == 8'hd8)? 32'h630c78ca
	         : (byte_in == 8'hd9)? 32'he9134912
	         : (byte_in == 8'hda)? 32'hf663df1c
	         : (byte_in == 8'hdb)? 32'h7c7ceec4
	         : (byte_in == 8'hdc)? 32'h7c1efcf9
	         : (byte_in == 8'hdd)? 32'hf601cd21
	         : (byte_in == 8'hde)? 32'he9715b2f
	         : (byte_in == 8'hdf)? 32'h636e6af7
	         : (byte_in == 8'he0)? 32'h5360ef7c
	         : (byte_in == 8'he1)? 32'hd97fdea4
	         : (byte_in == 8'he2)? 32'hc60f48aa
	         : (byte_in == 8'he3)? 32'h4c107972
	         : (byte_in == 8'he4)? 32'h4c726b4f
	         : (byte_in == 8'he5)? 32'hc66d5a97
	         : (byte_in == 8'he6)? 32'hd91dcc99
	         : (byte_in == 8'he7)? 32'h5302fd41
	         : (byte_in == 8'he8)? 32'h412b8742
	         : (byte_in == 8'he9)? 32'hcb34b69a
	         : (byte_in == 8'hea)? 32'hd4442094
	         : (byte_in == 8'heb)? 32'h5e5b114c
	         : (byte_in == 8'hec)? 32'h5e390371
	         : (byte_in == 8'hed)? 32'hd42632a9
	         : (byte_in == 8'hee)? 32'hcb56a4a7
	         : (byte_in == 8'hef)? 32'h4149957f
	         : (byte_in == 8'hf0)? 32'h5efd270b
	         : (byte_in == 8'hf1)? 32'hd4e216d3
	         : (byte_in == 8'hf2)? 32'hcb9280dd
	         : (byte_in == 8'hf3)? 32'h418db105
	         : (byte_in == 8'hf4)? 32'h41efa338
	         : (byte_in == 8'hf5)? 32'hcbf092e0
	         : (byte_in == 8'hf6)? 32'hd48004ee
	         : (byte_in == 8'hf7)? 32'h5e9f3536
	         : (byte_in == 8'hf8)? 32'h4cb64f35
	         : (byte_in == 8'hf9)? 32'hc6a97eed
	         : (byte_in == 8'hfa)? 32'hd9d9e8e3
	         : (byte_in == 8'hfb)? 32'h53c6d93b
	         : (byte_in == 8'hfc)? 32'h53a4cb06
	         : (byte_in == 8'hfd)? 32'hd9bbfade
	         : (byte_in == 8'hfe)? 32'hc6cb6cd0
	         :                     32'h4cd45d08;

endmodule
//}}}

module TABLE7(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h5a2b467e
	         : (byte_in == 8'h02)? 32'h90273769
	         : (byte_in == 8'h03)? 32'hca0c7117
	         : (byte_in == 8'h04)? 32'hb4578cfc
	         : (byte_in == 8'h05)? 32'hee7cca82
	         : (byte_in == 8'h06)? 32'h2470bb95
	         : (byte_in == 8'h07)? 32'h7e5bfdeb
	         : (byte_in == 8'h08)? 32'h204f6ed3
	         : (byte_in == 8'h09)? 32'h7a6428ad
	         : (byte_in == 8'h0a)? 32'hb06859ba
	         : (byte_in == 8'h0b)? 32'hea431fc4
	         : (byte_in == 8'h0c)? 32'h9418e22f
	         : (byte_in == 8'h0d)? 32'hce33a451
	         : (byte_in == 8'h0e)? 32'h043fd546
	         : (byte_in == 8'h0f)? 32'h5e149338
	         : (byte_in == 8'h10)? 32'h5b17d9e8
	         : (byte_in == 8'h11)? 32'h013c9f96
	         : (byte_in == 8'h12)? 32'hcb30ee81
	         : (byte_in == 8'h13)? 32'h911ba8ff
	         : (byte_in == 8'h14)? 32'hef405514
	         : (byte_in == 8'h15)? 32'hb56b136a
	         : (byte_in == 8'h16)? 32'h7f67627d
	         : (byte_in == 8'h17)? 32'h254c2403
	         : (byte_in == 8'h18)? 32'h7b58b73b
	         : (byte_in == 8'h19)? 32'h2173f145
	         : (byte_in == 8'h1a)? 32'heb7f8052
	         : (byte_in == 8'h1b)? 32'hb154c62c
	         : (byte_in == 8'h1c)? 32'hcf0f3bc7
	         : (byte_in == 8'h1d)? 32'h95247db9
	         : (byte_in == 8'h1e)? 32'h5f280cae
	         : (byte_in == 8'h1f)? 32'h05034ad0
	         : (byte_in == 8'h20)? 32'h4bb33a25
	         : (byte_in == 8'h21)? 32'h11987c5b
	         : (byte_in == 8'h22)? 32'hdb940d4c
	         : (byte_in == 8'h23)? 32'h81bf4b32
	         : (byte_in == 8'h24)? 32'hffe4b6d9
	         : (byte_in == 8'h25)? 32'ha5cff0a7
	         : (byte_in == 8'h26)? 32'h6fc381b0
	         : (byte_in == 8'h27)? 32'h35e8c7ce
	         : (byte_in == 8'h28)? 32'h6bfc54f6
	         : (byte_in == 8'h29)? 32'h31d71288
	         : (byte_in == 8'h2a)? 32'hfbdb639f
	         : (byte_in == 8'h2b)? 32'ha1f025e1
	         : (byte_in == 8'h2c)? 32'hdfabd80a
	         : (byte_in == 8'h2d)? 32'h85809e74
	         : (byte_in == 8'h2e)? 32'h4f8cef63
	         : (byte_in == 8'h2f)? 32'h15a7a91d
	         : (byte_in == 8'h30)? 32'h10a4e3cd
	         : (byte_in == 8'h31)? 32'h4a8fa5b3
	         : (byte_in == 8'h32)? 32'h8083d4a4
	         : (byte_in == 8'h33)? 32'hdaa892da
	         : (byte_in == 8'h34)? 32'ha4f36f31
	         : (byte_in == 8'h35)? 32'hfed8294f
	         : (byte_in == 8'h36)? 32'h34d45858
	         : (byte_in == 8'h37)? 32'h6eff1e26
	         : (byte_in == 8'h38)? 32'h30eb8d1e
	         : (byte_in == 8'h39)? 32'h6ac0cb60
	         : (byte_in == 8'h3a)? 32'ha0ccba77
	         : (byte_in == 8'h3b)? 32'hfae7fc09
	         : (byte_in == 8'h3c)? 32'h84bc01e2
	         : (byte_in == 8'h3d)? 32'hde97479c
	         : (byte_in == 8'h3e)? 32'h149b368b
	         : (byte_in == 8'h3f)? 32'h4eb070f5
	         : (byte_in == 8'h40)? 32'h859673c1
	         : (byte_in == 8'h41)? 32'hdfbd35bf
	         : (byte_in == 8'h42)? 32'h15b144a8
	         : (byte_in == 8'h43)? 32'h4f9a02d6
	         : (byte_in == 8'h44)? 32'h31c1ff3d
	         : (byte_in == 8'h45)? 32'h6beab943
	         : (byte_in == 8'h46)? 32'ha1e6c854
	         : (byte_in == 8'h47)? 32'hfbcd8e2a
	         : (byte_in == 8'h48)? 32'ha5d91d12
	         : (byte_in == 8'h49)? 32'hfff25b6c
	         : (byte_in == 8'h4a)? 32'h35fe2a7b
	         : (byte_in == 8'h4b)? 32'h6fd56c05
	         : (byte_in == 8'h4c)? 32'h118e91ee
	         : (byte_in == 8'h4d)? 32'h4ba5d790
	         : (byte_in == 8'h4e)? 32'h81a9a687
	         : (byte_in == 8'h4f)? 32'hdb82e0f9
	         : (byte_in == 8'h50)? 32'hde81aa29
	         : (byte_in == 8'h51)? 32'h84aaec57
	         : (byte_in == 8'h52)? 32'h4ea69d40
	         : (byte_in == 8'h53)? 32'h148ddb3e
	         : (byte_in == 8'h54)? 32'h6ad626d5
	         : (byte_in == 8'h55)? 32'h30fd60ab
	         : (byte_in == 8'h56)? 32'hfaf111bc
	         : (byte_in == 8'h57)? 32'ha0da57c2
	         : (byte_in == 8'h58)? 32'hfecec4fa
	         : (byte_in == 8'h59)? 32'ha4e58284
	         : (byte_in == 8'h5a)? 32'h6ee9f393
	         : (byte_in == 8'h5b)? 32'h34c2b5ed
	         : (byte_in == 8'h5c)? 32'h4a994806
	         : (byte_in == 8'h5d)? 32'h10b20e78
	         : (byte_in == 8'h5e)? 32'hdabe7f6f
	         : (byte_in == 8'h5f)? 32'h80953911
	         : (byte_in == 8'h60)? 32'hce2549e4
	         : (byte_in == 8'h61)? 32'h940e0f9a
	         : (byte_in == 8'h62)? 32'h5e027e8d
	         : (byte_in == 8'h63)? 32'h042938f3
	         : (byte_in == 8'h64)? 32'h7a72c518
	         : (byte_in == 8'h65)? 32'h20598366
	         : (byte_in == 8'h66)? 32'hea55f271
	         : (byte_in == 8'h67)? 32'hb07eb40f
	         : (byte_in == 8'h68)? 32'hee6a2737
	         : (byte_in == 8'h69)? 32'hb4416149
	         : (byte_in == 8'h6a)? 32'h7e4d105e
	         : (byte_in == 8'h6b)? 32'h24665620
	         : (byte_in == 8'h6c)? 32'h5a3dabcb
	         : (byte_in == 8'h6d)? 32'h0016edb5
	         : (byte_in == 8'h6e)? 32'hca1a9ca2
	         : (byte_in == 8'h6f)? 32'h9031dadc
	         : (byte_in == 8'h70)? 32'h9532900c
	         : (byte_in == 8'h71)? 32'hcf19d672
	         : (byte_in == 8'h72)? 32'h0515a765
	         : (byte_in == 8'h73)? 32'h5f3ee11b
	         : (byte_in == 8'h74)? 32'h21651cf0
	         : (byte_in == 8'h75)? 32'h7b4e5a8e
	         : (byte_in == 8'h76)? 32'hb1422b99
	         : (byte_in == 8'h77)? 32'heb696de7
	         : (byte_in == 8'h78)? 32'hb57dfedf
	         : (byte_in == 8'h79)? 32'hef56b8a1
	         : (byte_in == 8'h7a)? 32'h255ac9b6
	         : (byte_in == 8'h7b)? 32'h7f718fc8
	         : (byte_in == 8'h7c)? 32'h012a7223
	         : (byte_in == 8'h7d)? 32'h5b01345d
	         : (byte_in == 8'h7e)? 32'h910d454a
	         : (byte_in == 8'h7f)? 32'hcb260334
	         : (byte_in == 8'h80)? 32'h9c4a93c9
	         : (byte_in == 8'h81)? 32'hc661d5b7
	         : (byte_in == 8'h82)? 32'h0c6da4a0
	         : (byte_in == 8'h83)? 32'h5646e2de
	         : (byte_in == 8'h84)? 32'h281d1f35
	         : (byte_in == 8'h85)? 32'h7236594b
	         : (byte_in == 8'h86)? 32'hb83a285c
	         : (byte_in == 8'h87)? 32'he2116e22
	         : (byte_in == 8'h88)? 32'hbc05fd1a
	         : (byte_in == 8'h89)? 32'he62ebb64
	         : (byte_in == 8'h8a)? 32'h2c22ca73
	         : (byte_in == 8'h8b)? 32'h76098c0d
	         : (byte_in == 8'h8c)? 32'h085271e6
	         : (byte_in == 8'h8d)? 32'h52793798
	         : (byte_in == 8'h8e)? 32'h9875468f
	         : (byte_in == 8'h8f)? 32'hc25e00f1
	         : (byte_in == 8'h90)? 32'hc75d4a21
	         : (byte_in == 8'h91)? 32'h9d760c5f
	         : (byte_in == 8'h92)? 32'h577a7d48
	         : (byte_in == 8'h93)? 32'h0d513b36
	         : (byte_in == 8'h94)? 32'h730ac6dd
	         : (byte_in == 8'h95)? 32'h292180a3
	         : (byte_in == 8'h96)? 32'he32df1b4
	         : (byte_in == 8'h97)? 32'hb906b7ca
	         : (byte_in == 8'h98)? 32'he71224f2
	         : (byte_in == 8'h99)? 32'hbd39628c
	         : (byte_in == 8'h9a)? 32'h7735139b
	         : (byte_in == 8'h9b)? 32'h2d1e55e5
	         : (byte_in == 8'h9c)? 32'h5345a80e
	         : (byte_in == 8'h9d)? 32'h096eee70
	         : (byte_in == 8'h9e)? 32'hc3629f67
	         : (byte_in == 8'h9f)? 32'h9949d919
	         : (byte_in == 8'ha0)? 32'hd7f9a9ec
	         : (byte_in == 8'ha1)? 32'h8dd2ef92
	         : (byte_in == 8'ha2)? 32'h47de9e85
	         : (byte_in == 8'ha3)? 32'h1df5d8fb
	         : (byte_in == 8'ha4)? 32'h63ae2510
	         : (byte_in == 8'ha5)? 32'h3985636e
	         : (byte_in == 8'ha6)? 32'hf3891279
	         : (byte_in == 8'ha7)? 32'ha9a25407
	         : (byte_in == 8'ha8)? 32'hf7b6c73f
	         : (byte_in == 8'ha9)? 32'had9d8141
	         : (byte_in == 8'haa)? 32'h6791f056
	         : (byte_in == 8'hab)? 32'h3dbab628
	         : (byte_in == 8'hac)? 32'h43e14bc3
	         : (byte_in == 8'had)? 32'h19ca0dbd
	         : (byte_in == 8'hae)? 32'hd3c67caa
	         : (byte_in == 8'haf)? 32'h89ed3ad4
	         : (byte_in == 8'hb0)? 32'h8cee7004
	         : (byte_in == 8'hb1)? 32'hd6c5367a
	         : (byte_in == 8'hb2)? 32'h1cc9476d
	         : (byte_in == 8'hb3)? 32'h46e20113
	         : (byte_in == 8'hb4)? 32'h38b9fcf8
	         : (byte_in == 8'hb5)? 32'h6292ba86
	         : (byte_in == 8'hb6)? 32'ha89ecb91
	         : (byte_in == 8'hb7)? 32'hf2b58def
	         : (byte_in == 8'hb8)? 32'haca11ed7
	         : (byte_in == 8'hb9)? 32'hf68a58a9
	         : (byte_in == 8'hba)? 32'h3c8629be
	         : (byte_in == 8'hbb)? 32'h66ad6fc0
	         : (byte_in == 8'hbc)? 32'h18f6922b
	         : (byte_in == 8'hbd)? 32'h42ddd455
	         : (byte_in == 8'hbe)? 32'h88d1a542
	         : (byte_in == 8'hbf)? 32'hd2fae33c
	         : (byte_in == 8'hc0)? 32'h19dce008
	         : (byte_in == 8'hc1)? 32'h43f7a676
	         : (byte_in == 8'hc2)? 32'h89fbd761
	         : (byte_in == 8'hc3)? 32'hd3d0911f
	         : (byte_in == 8'hc4)? 32'had8b6cf4
	         : (byte_in == 8'hc5)? 32'hf7a02a8a
	         : (byte_in == 8'hc6)? 32'h3dac5b9d
	         : (byte_in == 8'hc7)? 32'h67871de3
	         : (byte_in == 8'hc8)? 32'h39938edb
	         : (byte_in == 8'hc9)? 32'h63b8c8a5
	         : (byte_in == 8'hca)? 32'ha9b4b9b2
	         : (byte_in == 8'hcb)? 32'hf39fffcc
	         : (byte_in == 8'hcc)? 32'h8dc40227
	         : (byte_in == 8'hcd)? 32'hd7ef4459
	         : (byte_in == 8'hce)? 32'h1de3354e
	         : (byte_in == 8'hcf)? 32'h47c87330
	         : (byte_in == 8'hd0)? 32'h42cb39e0
	         : (byte_in == 8'hd1)? 32'h18e07f9e
	         : (byte_in == 8'hd2)? 32'hd2ec0e89
	         : (byte_in == 8'hd3)? 32'h88c748f7
	         : (byte_in == 8'hd4)? 32'hf69cb51c
	         : (byte_in == 8'hd5)? 32'hacb7f362
	         : (byte_in == 8'hd6)? 32'h66bb8275
	         : (byte_in == 8'hd7)? 32'h3c90c40b
	         : (byte_in == 8'hd8)? 32'h62845733
	         : (byte_in == 8'hd9)? 32'h38af114d
	         : (byte_in == 8'hda)? 32'hf2a3605a
	         : (byte_in == 8'hdb)? 32'ha8882624
	         : (byte_in == 8'hdc)? 32'hd6d3dbcf
	         : (byte_in == 8'hdd)? 32'h8cf89db1
	         : (byte_in == 8'hde)? 32'h46f4eca6
	         : (byte_in == 8'hdf)? 32'h1cdfaad8
	         : (byte_in == 8'he0)? 32'h526fda2d
	         : (byte_in == 8'he1)? 32'h08449c53
	         : (byte_in == 8'he2)? 32'hc248ed44
	         : (byte_in == 8'he3)? 32'h9863ab3a
	         : (byte_in == 8'he4)? 32'he63856d1
	         : (byte_in == 8'he5)? 32'hbc1310af
	         : (byte_in == 8'he6)? 32'h761f61b8
	         : (byte_in == 8'he7)? 32'h2c3427c6
	         : (byte_in == 8'he8)? 32'h7220b4fe
	         : (byte_in == 8'he9)? 32'h280bf280
	         : (byte_in == 8'hea)? 32'he2078397
	         : (byte_in == 8'heb)? 32'hb82cc5e9
	         : (byte_in == 8'hec)? 32'hc6773802
	         : (byte_in == 8'hed)? 32'h9c5c7e7c
	         : (byte_in == 8'hee)? 32'h56500f6b
	         : (byte_in == 8'hef)? 32'h0c7b4915
	         : (byte_in == 8'hf0)? 32'h097803c5
	         : (byte_in == 8'hf1)? 32'h535345bb
	         : (byte_in == 8'hf2)? 32'h995f34ac
	         : (byte_in == 8'hf3)? 32'hc37472d2
	         : (byte_in == 8'hf4)? 32'hbd2f8f39
	         : (byte_in == 8'hf5)? 32'he704c947
	         : (byte_in == 8'hf6)? 32'h2d08b850
	         : (byte_in == 8'hf7)? 32'h7723fe2e
	         : (byte_in == 8'hf8)? 32'h29376d16
	         : (byte_in == 8'hf9)? 32'h731c2b68
	         : (byte_in == 8'hfa)? 32'hb9105a7f
	         : (byte_in == 8'hfb)? 32'he33b1c01
	         : (byte_in == 8'hfc)? 32'h9d60e1ea
	         : (byte_in == 8'hfd)? 32'hc74ba794
	         : (byte_in == 8'hfe)? 32'h0d47d683
	         :                     32'h576c90fd;

endmodule
//}}}

module TABLE8(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'hae0ebb05
	         : (byte_in == 8'h02)? 32'h6bf648a4
	         : (byte_in == 8'h03)? 32'hc5f8f3a1
	         : (byte_in == 8'h04)? 32'h99e585aa
	         : (byte_in == 8'h05)? 32'h37eb3eaf
	         : (byte_in == 8'h06)? 32'hf213cd0e
	         : (byte_in == 8'h07)? 32'h5c1d760b
	         : (byte_in == 8'h08)? 32'h79e22a4c
	         : (byte_in == 8'h09)? 32'hd7ec9149
	         : (byte_in == 8'h0a)? 32'h121462e8
	         : (byte_in == 8'h0b)? 32'hbc1ad9ed
	         : (byte_in == 8'h0c)? 32'he007afe6
	         : (byte_in == 8'h0d)? 32'h4e0914e3
	         : (byte_in == 8'h0e)? 32'h8bf1e742
	         : (byte_in == 8'h0f)? 32'h25ff5c47
	         : (byte_in == 8'h10)? 32'h9dc5b050
	         : (byte_in == 8'h11)? 32'h33cb0b55
	         : (byte_in == 8'h12)? 32'hf633f8f4
	         : (byte_in == 8'h13)? 32'h583d43f1
	         : (byte_in == 8'h14)? 32'h042035fa
	         : (byte_in == 8'h15)? 32'haa2e8eff
	         : (byte_in == 8'h16)? 32'h6fd67d5e
	         : (byte_in == 8'h17)? 32'hc1d8c65b
	         : (byte_in == 8'h18)? 32'he4279a1c
	         : (byte_in == 8'h19)? 32'h4a292119
	         : (byte_in == 8'h1a)? 32'h8fd1d2b8
	         : (byte_in == 8'h1b)? 32'h21df69bd
	         : (byte_in == 8'h1c)? 32'h7dc21fb6
	         : (byte_in == 8'h1d)? 32'hd3cca4b3
	         : (byte_in == 8'h1e)? 32'h16345712
	         : (byte_in == 8'h1f)? 32'hb83aec17
	         : (byte_in == 8'h20)? 32'h98321c3d
	         : (byte_in == 8'h21)? 32'h363ca738
	         : (byte_in == 8'h22)? 32'hf3c45499
	         : (byte_in == 8'h23)? 32'h5dcaef9c
	         : (byte_in == 8'h24)? 32'h01d79997
	         : (byte_in == 8'h25)? 32'hafd92292
	         : (byte_in == 8'h26)? 32'h6a21d133
	         : (byte_in == 8'h27)? 32'hc42f6a36
	         : (byte_in == 8'h28)? 32'he1d03671
	         : (byte_in == 8'h29)? 32'h4fde8d74
	         : (byte_in == 8'h2a)? 32'h8a267ed5
	         : (byte_in == 8'h2b)? 32'h2428c5d0
	         : (byte_in == 8'h2c)? 32'h7835b3db
	         : (byte_in == 8'h2d)? 32'hd63b08de
	         : (byte_in == 8'h2e)? 32'h13c3fb7f
	         : (byte_in == 8'h2f)? 32'hbdcd407a
	         : (byte_in == 8'h30)? 32'h05f7ac6d
	         : (byte_in == 8'h31)? 32'habf91768
	         : (byte_in == 8'h32)? 32'h6e01e4c9
	         : (byte_in == 8'h33)? 32'hc00f5fcc
	         : (byte_in == 8'h34)? 32'h9c1229c7
	         : (byte_in == 8'h35)? 32'h321c92c2
	         : (byte_in == 8'h36)? 32'hf7e46163
	         : (byte_in == 8'h37)? 32'h59eada66
	         : (byte_in == 8'h38)? 32'h7c158621
	         : (byte_in == 8'h39)? 32'hd21b3d24
	         : (byte_in == 8'h3a)? 32'h17e3ce85
	         : (byte_in == 8'h3b)? 32'hb9ed7580
	         : (byte_in == 8'h3c)? 32'he5f0038b
	         : (byte_in == 8'h3d)? 32'h4bfeb88e
	         : (byte_in == 8'h3e)? 32'h8e064b2f
	         : (byte_in == 8'h3f)? 32'h2008f02a
	         : (byte_in == 8'h40)? 32'hfe739301
	         : (byte_in == 8'h41)? 32'h507d2804
	         : (byte_in == 8'h42)? 32'h9585dba5
	         : (byte_in == 8'h43)? 32'h3b8b60a0
	         : (byte_in == 8'h44)? 32'h679616ab
	         : (byte_in == 8'h45)? 32'hc998adae
	         : (byte_in == 8'h46)? 32'h0c605e0f
	         : (byte_in == 8'h47)? 32'ha26ee50a
	         : (byte_in == 8'h48)? 32'h8791b94d
	         : (byte_in == 8'h49)? 32'h299f0248
	         : (byte_in == 8'h4a)? 32'hec67f1e9
	         : (byte_in == 8'h4b)? 32'h42694aec
	         : (byte_in == 8'h4c)? 32'h1e743ce7
	         : (byte_in == 8'h4d)? 32'hb07a87e2
	         : (byte_in == 8'h4e)? 32'h75827443
	         : (byte_in == 8'h4f)? 32'hdb8ccf46
	         : (byte_in == 8'h50)? 32'h63b62351
	         : (byte_in == 8'h51)? 32'hcdb89854
	         : (byte_in == 8'h52)? 32'h08406bf5
	         : (byte_in == 8'h53)? 32'ha64ed0f0
	         : (byte_in == 8'h54)? 32'hfa53a6fb
	         : (byte_in == 8'h55)? 32'h545d1dfe
	         : (byte_in == 8'h56)? 32'h91a5ee5f
	         : (byte_in == 8'h57)? 32'h3fab555a
	         : (byte_in == 8'h58)? 32'h1a54091d
	         : (byte_in == 8'h59)? 32'hb45ab218
	         : (byte_in == 8'h5a)? 32'h71a241b9
	         : (byte_in == 8'h5b)? 32'hdfacfabc
	         : (byte_in == 8'h5c)? 32'h83b18cb7
	         : (byte_in == 8'h5d)? 32'h2dbf37b2
	         : (byte_in == 8'h5e)? 32'he847c413
	         : (byte_in == 8'h5f)? 32'h46497f16
	         : (byte_in == 8'h60)? 32'h66418f3c
	         : (byte_in == 8'h61)? 32'hc84f3439
	         : (byte_in == 8'h62)? 32'h0db7c798
	         : (byte_in == 8'h63)? 32'ha3b97c9d
	         : (byte_in == 8'h64)? 32'hffa40a96
	         : (byte_in == 8'h65)? 32'h51aab193
	         : (byte_in == 8'h66)? 32'h94524232
	         : (byte_in == 8'h67)? 32'h3a5cf937
	         : (byte_in == 8'h68)? 32'h1fa3a570
	         : (byte_in == 8'h69)? 32'hb1ad1e75
	         : (byte_in == 8'h6a)? 32'h7455edd4
	         : (byte_in == 8'h6b)? 32'hda5b56d1
	         : (byte_in == 8'h6c)? 32'h864620da
	         : (byte_in == 8'h6d)? 32'h28489bdf
	         : (byte_in == 8'h6e)? 32'hedb0687e
	         : (byte_in == 8'h6f)? 32'h43bed37b
	         : (byte_in == 8'h70)? 32'hfb843f6c
	         : (byte_in == 8'h71)? 32'h558a8469
	         : (byte_in == 8'h72)? 32'h907277c8
	         : (byte_in == 8'h73)? 32'h3e7ccccd
	         : (byte_in == 8'h74)? 32'h6261bac6
	         : (byte_in == 8'h75)? 32'hcc6f01c3
	         : (byte_in == 8'h76)? 32'h0997f262
	         : (byte_in == 8'h77)? 32'ha7994967
	         : (byte_in == 8'h78)? 32'h82661520
	         : (byte_in == 8'h79)? 32'h2c68ae25
	         : (byte_in == 8'h7a)? 32'he9905d84
	         : (byte_in == 8'h7b)? 32'h479ee681
	         : (byte_in == 8'h7c)? 32'h1b83908a
	         : (byte_in == 8'h7d)? 32'hb58d2b8f
	         : (byte_in == 8'h7e)? 32'h7075d82e
	         : (byte_in == 8'h7f)? 32'hde7b632b
	         : (byte_in == 8'h80)? 32'h9e6a837e
	         : (byte_in == 8'h81)? 32'h3064387b
	         : (byte_in == 8'h82)? 32'hf59ccbda
	         : (byte_in == 8'h83)? 32'h5b9270df
	         : (byte_in == 8'h84)? 32'h078f06d4
	         : (byte_in == 8'h85)? 32'ha981bdd1
	         : (byte_in == 8'h86)? 32'h6c794e70
	         : (byte_in == 8'h87)? 32'hc277f575
	         : (byte_in == 8'h88)? 32'he788a932
	         : (byte_in == 8'h89)? 32'h49861237
	         : (byte_in == 8'h8a)? 32'h8c7ee196
	         : (byte_in == 8'h8b)? 32'h22705a93
	         : (byte_in == 8'h8c)? 32'h7e6d2c98
	         : (byte_in == 8'h8d)? 32'hd063979d
	         : (byte_in == 8'h8e)? 32'h159b643c
	         : (byte_in == 8'h8f)? 32'hbb95df39
	         : (byte_in == 8'h90)? 32'h03af332e
	         : (byte_in == 8'h91)? 32'hada1882b
	         : (byte_in == 8'h92)? 32'h68597b8a
	         : (byte_in == 8'h93)? 32'hc657c08f
	         : (byte_in == 8'h94)? 32'h9a4ab684
	         : (byte_in == 8'h95)? 32'h34440d81
	         : (byte_in == 8'h96)? 32'hf1bcfe20
	         : (byte_in == 8'h97)? 32'h5fb24525
	         : (byte_in == 8'h98)? 32'h7a4d1962
	         : (byte_in == 8'h99)? 32'hd443a267
	         : (byte_in == 8'h9a)? 32'h11bb51c6
	         : (byte_in == 8'h9b)? 32'hbfb5eac3
	         : (byte_in == 8'h9c)? 32'he3a89cc8
	         : (byte_in == 8'h9d)? 32'h4da627cd
	         : (byte_in == 8'h9e)? 32'h885ed46c
	         : (byte_in == 8'h9f)? 32'h26506f69
	         : (byte_in == 8'ha0)? 32'h06589f43
	         : (byte_in == 8'ha1)? 32'ha8562446
	         : (byte_in == 8'ha2)? 32'h6daed7e7
	         : (byte_in == 8'ha3)? 32'hc3a06ce2
	         : (byte_in == 8'ha4)? 32'h9fbd1ae9
	         : (byte_in == 8'ha5)? 32'h31b3a1ec
	         : (byte_in == 8'ha6)? 32'hf44b524d
	         : (byte_in == 8'ha7)? 32'h5a45e948
	         : (byte_in == 8'ha8)? 32'h7fbab50f
	         : (byte_in == 8'ha9)? 32'hd1b40e0a
	         : (byte_in == 8'haa)? 32'h144cfdab
	         : (byte_in == 8'hab)? 32'hba4246ae
	         : (byte_in == 8'hac)? 32'he65f30a5
	         : (byte_in == 8'had)? 32'h48518ba0
	         : (byte_in == 8'hae)? 32'h8da97801
	         : (byte_in == 8'haf)? 32'h23a7c304
	         : (byte_in == 8'hb0)? 32'h9b9d2f13
	         : (byte_in == 8'hb1)? 32'h35939416
	         : (byte_in == 8'hb2)? 32'hf06b67b7
	         : (byte_in == 8'hb3)? 32'h5e65dcb2
	         : (byte_in == 8'hb4)? 32'h0278aab9
	         : (byte_in == 8'hb5)? 32'hac7611bc
	         : (byte_in == 8'hb6)? 32'h698ee21d
	         : (byte_in == 8'hb7)? 32'hc7805918
	         : (byte_in == 8'hb8)? 32'he27f055f
	         : (byte_in == 8'hb9)? 32'h4c71be5a
	         : (byte_in == 8'hba)? 32'h89894dfb
	         : (byte_in == 8'hbb)? 32'h2787f6fe
	         : (byte_in == 8'hbc)? 32'h7b9a80f5
	         : (byte_in == 8'hbd)? 32'hd5943bf0
	         : (byte_in == 8'hbe)? 32'h106cc851
	         : (byte_in == 8'hbf)? 32'hbe627354
	         : (byte_in == 8'hc0)? 32'h6019107f
	         : (byte_in == 8'hc1)? 32'hce17ab7a
	         : (byte_in == 8'hc2)? 32'h0bef58db
	         : (byte_in == 8'hc3)? 32'ha5e1e3de
	         : (byte_in == 8'hc4)? 32'hf9fc95d5
	         : (byte_in == 8'hc5)? 32'h57f22ed0
	         : (byte_in == 8'hc6)? 32'h920add71
	         : (byte_in == 8'hc7)? 32'h3c046674
	         : (byte_in == 8'hc8)? 32'h19fb3a33
	         : (byte_in == 8'hc9)? 32'hb7f58136
	         : (byte_in == 8'hca)? 32'h720d7297
	         : (byte_in == 8'hcb)? 32'hdc03c992
	         : (byte_in == 8'hcc)? 32'h801ebf99
	         : (byte_in == 8'hcd)? 32'h2e10049c
	         : (byte_in == 8'hce)? 32'hebe8f73d
	         : (byte_in == 8'hcf)? 32'h45e64c38
	         : (byte_in == 8'hd0)? 32'hfddca02f
	         : (byte_in == 8'hd1)? 32'h53d21b2a
	         : (byte_in == 8'hd2)? 32'h962ae88b
	         : (byte_in == 8'hd3)? 32'h3824538e
	         : (byte_in == 8'hd4)? 32'h64392585
	         : (byte_in == 8'hd5)? 32'hca379e80
	         : (byte_in == 8'hd6)? 32'h0fcf6d21
	         : (byte_in == 8'hd7)? 32'ha1c1d624
	         : (byte_in == 8'hd8)? 32'h843e8a63
	         : (byte_in == 8'hd9)? 32'h2a303166
	         : (byte_in == 8'hda)? 32'hefc8c2c7
	         : (byte_in == 8'hdb)? 32'h41c679c2
	         : (byte_in == 8'hdc)? 32'h1ddb0fc9
	         : (byte_in == 8'hdd)? 32'hb3d5b4cc
	         : (byte_in == 8'hde)? 32'h762d476d
	         : (byte_in == 8'hdf)? 32'hd823fc68
	         : (byte_in == 8'he0)? 32'hf82b0c42
	         : (byte_in == 8'he1)? 32'h5625b747
	         : (byte_in == 8'he2)? 32'h93dd44e6
	         : (byte_in == 8'he3)? 32'h3dd3ffe3
	         : (byte_in == 8'he4)? 32'h61ce89e8
	         : (byte_in == 8'he5)? 32'hcfc032ed
	         : (byte_in == 8'he6)? 32'h0a38c14c
	         : (byte_in == 8'he7)? 32'ha4367a49
	         : (byte_in == 8'he8)? 32'h81c9260e
	         : (byte_in == 8'he9)? 32'h2fc79d0b
	         : (byte_in == 8'hea)? 32'hea3f6eaa
	         : (byte_in == 8'heb)? 32'h4431d5af
	         : (byte_in == 8'hec)? 32'h182ca3a4
	         : (byte_in == 8'hed)? 32'hb62218a1
	         : (byte_in == 8'hee)? 32'h73daeb00
	         : (byte_in == 8'hef)? 32'hddd45005
	         : (byte_in == 8'hf0)? 32'h65eebc12
	         : (byte_in == 8'hf1)? 32'hcbe00717
	         : (byte_in == 8'hf2)? 32'h0e18f4b6
	         : (byte_in == 8'hf3)? 32'ha0164fb3
	         : (byte_in == 8'hf4)? 32'hfc0b39b8
	         : (byte_in == 8'hf5)? 32'h520582bd
	         : (byte_in == 8'hf6)? 32'h97fd711c
	         : (byte_in == 8'hf7)? 32'h39f3ca19
	         : (byte_in == 8'hf8)? 32'h1c0c965e
	         : (byte_in == 8'hf9)? 32'hb2022d5b
	         : (byte_in == 8'hfa)? 32'h77fadefa
	         : (byte_in == 8'hfb)? 32'hd9f465ff
	         : (byte_in == 8'hfc)? 32'h85e913f4
	         : (byte_in == 8'hfd)? 32'h2be7a8f1
	         : (byte_in == 8'hfe)? 32'hee1f5b50
	         :                     32'h4011e055;

endmodule
//}}}

module TABLE9(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'hfce72602
	         : (byte_in == 8'h02)? 32'h3cd406fc
	         : (byte_in == 8'h03)? 32'hc03320fe
	         : (byte_in == 8'h04)? 32'hf9ce4c04
	         : (byte_in == 8'h05)? 32'h05296a06
	         : (byte_in == 8'h06)? 32'hc51a4af8
	         : (byte_in == 8'h07)? 32'h39fd6cfa
	         : (byte_in == 8'h08)? 32'h79a90df9
	         : (byte_in == 8'h09)? 32'h854e2bfb
	         : (byte_in == 8'h0a)? 32'h457d0b05
	         : (byte_in == 8'h0b)? 32'hb99a2d07
	         : (byte_in == 8'h0c)? 32'h806741fd
	         : (byte_in == 8'h0d)? 32'h7c8067ff
	         : (byte_in == 8'h0e)? 32'hbcb34701
	         : (byte_in == 8'h0f)? 32'h40546103
	         : (byte_in == 8'h10)? 32'h36656ba8
	         : (byte_in == 8'h11)? 32'hca824daa
	         : (byte_in == 8'h12)? 32'h0ab16d54
	         : (byte_in == 8'h13)? 32'hf6564b56
	         : (byte_in == 8'h14)? 32'hcfab27ac
	         : (byte_in == 8'h15)? 32'h334c01ae
	         : (byte_in == 8'h16)? 32'hf37f2150
	         : (byte_in == 8'h17)? 32'h0f980752
	         : (byte_in == 8'h18)? 32'h4fcc6651
	         : (byte_in == 8'h19)? 32'hb32b4053
	         : (byte_in == 8'h1a)? 32'h731860ad
	         : (byte_in == 8'h1b)? 32'h8fff46af
	         : (byte_in == 8'h1c)? 32'hb6022a55
	         : (byte_in == 8'h1d)? 32'h4ae50c57
	         : (byte_in == 8'h1e)? 32'h8ad62ca9
	         : (byte_in == 8'h1f)? 32'h76310aab
	         : (byte_in == 8'h20)? 32'h5d5ca0f7
	         : (byte_in == 8'h21)? 32'ha1bb86f5
	         : (byte_in == 8'h22)? 32'h6188a60b
	         : (byte_in == 8'h23)? 32'h9d6f8009
	         : (byte_in == 8'h24)? 32'ha492ecf3
	         : (byte_in == 8'h25)? 32'h5875caf1
	         : (byte_in == 8'h26)? 32'h9846ea0f
	         : (byte_in == 8'h27)? 32'h64a1cc0d
	         : (byte_in == 8'h28)? 32'h24f5ad0e
	         : (byte_in == 8'h29)? 32'hd8128b0c
	         : (byte_in == 8'h2a)? 32'h1821abf2
	         : (byte_in == 8'h2b)? 32'he4c68df0
	         : (byte_in == 8'h2c)? 32'hdd3be10a
	         : (byte_in == 8'h2d)? 32'h21dcc708
	         : (byte_in == 8'h2e)? 32'he1efe7f6
	         : (byte_in == 8'h2f)? 32'h1d08c1f4
	         : (byte_in == 8'h30)? 32'h6b39cb5f
	         : (byte_in == 8'h31)? 32'h97deed5d
	         : (byte_in == 8'h32)? 32'h57edcda3
	         : (byte_in == 8'h33)? 32'hab0aeba1
	         : (byte_in == 8'h34)? 32'h92f7875b
	         : (byte_in == 8'h35)? 32'h6e10a159
	         : (byte_in == 8'h36)? 32'hae2381a7
	         : (byte_in == 8'h37)? 32'h52c4a7a5
	         : (byte_in == 8'h38)? 32'h1290c6a6
	         : (byte_in == 8'h39)? 32'hee77e0a4
	         : (byte_in == 8'h3a)? 32'h2e44c05a
	         : (byte_in == 8'h3b)? 32'hd2a3e658
	         : (byte_in == 8'h3c)? 32'heb5e8aa2
	         : (byte_in == 8'h3d)? 32'h17b9aca0
	         : (byte_in == 8'h3e)? 32'hd78a8c5e
	         : (byte_in == 8'h3f)? 32'h2b6daa5c
	         : (byte_in == 8'h40)? 32'hc2c46c55
	         : (byte_in == 8'h41)? 32'h3e234a57
	         : (byte_in == 8'h42)? 32'hfe106aa9
	         : (byte_in == 8'h43)? 32'h02f74cab
	         : (byte_in == 8'h44)? 32'h3b0a2051
	         : (byte_in == 8'h45)? 32'hc7ed0653
	         : (byte_in == 8'h46)? 32'h07de26ad
	         : (byte_in == 8'h47)? 32'hfb3900af
	         : (byte_in == 8'h48)? 32'hbb6d61ac
	         : (byte_in == 8'h49)? 32'h478a47ae
	         : (byte_in == 8'h4a)? 32'h87b96750
	         : (byte_in == 8'h4b)? 32'h7b5e4152
	         : (byte_in == 8'h4c)? 32'h42a32da8
	         : (byte_in == 8'h4d)? 32'hbe440baa
	         : (byte_in == 8'h4e)? 32'h7e772b54
	         : (byte_in == 8'h4f)? 32'h82900d56
	         : (byte_in == 8'h50)? 32'hf4a107fd
	         : (byte_in == 8'h51)? 32'h084621ff
	         : (byte_in == 8'h52)? 32'hc8750101
	         : (byte_in == 8'h53)? 32'h34922703
	         : (byte_in == 8'h54)? 32'h0d6f4bf9
	         : (byte_in == 8'h55)? 32'hf1886dfb
	         : (byte_in == 8'h56)? 32'h31bb4d05
	         : (byte_in == 8'h57)? 32'hcd5c6b07
	         : (byte_in == 8'h58)? 32'h8d080a04
	         : (byte_in == 8'h59)? 32'h71ef2c06
	         : (byte_in == 8'h5a)? 32'hb1dc0cf8
	         : (byte_in == 8'h5b)? 32'h4d3b2afa
	         : (byte_in == 8'h5c)? 32'h74c64600
	         : (byte_in == 8'h5d)? 32'h88216002
	         : (byte_in == 8'h5e)? 32'h481240fc
	         : (byte_in == 8'h5f)? 32'hb4f566fe
	         : (byte_in == 8'h60)? 32'h9f98cca2
	         : (byte_in == 8'h61)? 32'h637feaa0
	         : (byte_in == 8'h62)? 32'ha34cca5e
	         : (byte_in == 8'h63)? 32'h5fabec5c
	         : (byte_in == 8'h64)? 32'h665680a6
	         : (byte_in == 8'h65)? 32'h9ab1a6a4
	         : (byte_in == 8'h66)? 32'h5a82865a
	         : (byte_in == 8'h67)? 32'ha665a058
	         : (byte_in == 8'h68)? 32'he631c15b
	         : (byte_in == 8'h69)? 32'h1ad6e759
	         : (byte_in == 8'h6a)? 32'hdae5c7a7
	         : (byte_in == 8'h6b)? 32'h2602e1a5
	         : (byte_in == 8'h6c)? 32'h1fff8d5f
	         : (byte_in == 8'h6d)? 32'he318ab5d
	         : (byte_in == 8'h6e)? 32'h232b8ba3
	         : (byte_in == 8'h6f)? 32'hdfccada1
	         : (byte_in == 8'h70)? 32'ha9fda70a
	         : (byte_in == 8'h71)? 32'h551a8108
	         : (byte_in == 8'h72)? 32'h9529a1f6
	         : (byte_in == 8'h73)? 32'h69ce87f4
	         : (byte_in == 8'h74)? 32'h5033eb0e
	         : (byte_in == 8'h75)? 32'hacd4cd0c
	         : (byte_in == 8'h76)? 32'h6ce7edf2
	         : (byte_in == 8'h77)? 32'h9000cbf0
	         : (byte_in == 8'h78)? 32'hd054aaf3
	         : (byte_in == 8'h79)? 32'h2cb38cf1
	         : (byte_in == 8'h7a)? 32'hec80ac0f
	         : (byte_in == 8'h7b)? 32'h10678a0d
	         : (byte_in == 8'h7c)? 32'h299ae6f7
	         : (byte_in == 8'h7d)? 32'hd57dc0f5
	         : (byte_in == 8'h7e)? 32'h154ee00b
	         : (byte_in == 8'h7f)? 32'he9a9c609
	         : (byte_in == 8'h80)? 32'hd14e094b
	         : (byte_in == 8'h81)? 32'h2da92f49
	         : (byte_in == 8'h82)? 32'hed9a0fb7
	         : (byte_in == 8'h83)? 32'h117d29b5
	         : (byte_in == 8'h84)? 32'h2880454f
	         : (byte_in == 8'h85)? 32'hd467634d
	         : (byte_in == 8'h86)? 32'h145443b3
	         : (byte_in == 8'h87)? 32'he8b365b1
	         : (byte_in == 8'h88)? 32'ha8e704b2
	         : (byte_in == 8'h89)? 32'h540022b0
	         : (byte_in == 8'h8a)? 32'h9433024e
	         : (byte_in == 8'h8b)? 32'h68d4244c
	         : (byte_in == 8'h8c)? 32'h512948b6
	         : (byte_in == 8'h8d)? 32'hadce6eb4
	         : (byte_in == 8'h8e)? 32'h6dfd4e4a
	         : (byte_in == 8'h8f)? 32'h911a6848
	         : (byte_in == 8'h90)? 32'he72b62e3
	         : (byte_in == 8'h91)? 32'h1bcc44e1
	         : (byte_in == 8'h92)? 32'hdbff641f
	         : (byte_in == 8'h93)? 32'h2718421d
	         : (byte_in == 8'h94)? 32'h1ee52ee7
	         : (byte_in == 8'h95)? 32'he20208e5
	         : (byte_in == 8'h96)? 32'h2231281b
	         : (byte_in == 8'h97)? 32'hded60e19
	         : (byte_in == 8'h98)? 32'h9e826f1a
	         : (byte_in == 8'h99)? 32'h62654918
	         : (byte_in == 8'h9a)? 32'ha25669e6
	         : (byte_in == 8'h9b)? 32'h5eb14fe4
	         : (byte_in == 8'h9c)? 32'h674c231e
	         : (byte_in == 8'h9d)? 32'h9bab051c
	         : (byte_in == 8'h9e)? 32'h5b9825e2
	         : (byte_in == 8'h9f)? 32'ha77f03e0
	         : (byte_in == 8'ha0)? 32'h8c12a9bc
	         : (byte_in == 8'ha1)? 32'h70f58fbe
	         : (byte_in == 8'ha2)? 32'hb0c6af40
	         : (byte_in == 8'ha3)? 32'h4c218942
	         : (byte_in == 8'ha4)? 32'h75dce5b8
	         : (byte_in == 8'ha5)? 32'h893bc3ba
	         : (byte_in == 8'ha6)? 32'h4908e344
	         : (byte_in == 8'ha7)? 32'hb5efc546
	         : (byte_in == 8'ha8)? 32'hf5bba445
	         : (byte_in == 8'ha9)? 32'h095c8247
	         : (byte_in == 8'haa)? 32'hc96fa2b9
	         : (byte_in == 8'hab)? 32'h358884bb
	         : (byte_in == 8'hac)? 32'h0c75e841
	         : (byte_in == 8'had)? 32'hf092ce43
	         : (byte_in == 8'hae)? 32'h30a1eebd
	         : (byte_in == 8'haf)? 32'hcc46c8bf
	         : (byte_in == 8'hb0)? 32'hba77c214
	         : (byte_in == 8'hb1)? 32'h4690e416
	         : (byte_in == 8'hb2)? 32'h86a3c4e8
	         : (byte_in == 8'hb3)? 32'h7a44e2ea
	         : (byte_in == 8'hb4)? 32'h43b98e10
	         : (byte_in == 8'hb5)? 32'hbf5ea812
	         : (byte_in == 8'hb6)? 32'h7f6d88ec
	         : (byte_in == 8'hb7)? 32'h838aaeee
	         : (byte_in == 8'hb8)? 32'hc3decfed
	         : (byte_in == 8'hb9)? 32'h3f39e9ef
	         : (byte_in == 8'hba)? 32'hff0ac911
	         : (byte_in == 8'hbb)? 32'h03edef13
	         : (byte_in == 8'hbc)? 32'h3a1083e9
	         : (byte_in == 8'hbd)? 32'hc6f7a5eb
	         : (byte_in == 8'hbe)? 32'h06c48515
	         : (byte_in == 8'hbf)? 32'hfa23a317
	         : (byte_in == 8'hc0)? 32'h138a651e
	         : (byte_in == 8'hc1)? 32'hef6d431c
	         : (byte_in == 8'hc2)? 32'h2f5e63e2
	         : (byte_in == 8'hc3)? 32'hd3b945e0
	         : (byte_in == 8'hc4)? 32'hea44291a
	         : (byte_in == 8'hc5)? 32'h16a30f18
	         : (byte_in == 8'hc6)? 32'hd6902fe6
	         : (byte_in == 8'hc7)? 32'h2a7709e4
	         : (byte_in == 8'hc8)? 32'h6a2368e7
	         : (byte_in == 8'hc9)? 32'h96c44ee5
	         : (byte_in == 8'hca)? 32'h56f76e1b
	         : (byte_in == 8'hcb)? 32'haa104819
	         : (byte_in == 8'hcc)? 32'h93ed24e3
	         : (byte_in == 8'hcd)? 32'h6f0a02e1
	         : (byte_in == 8'hce)? 32'haf39221f
	         : (byte_in == 8'hcf)? 32'h53de041d
	         : (byte_in == 8'hd0)? 32'h25ef0eb6
	         : (byte_in == 8'hd1)? 32'hd90828b4
	         : (byte_in == 8'hd2)? 32'h193b084a
	         : (byte_in == 8'hd3)? 32'he5dc2e48
	         : (byte_in == 8'hd4)? 32'hdc2142b2
	         : (byte_in == 8'hd5)? 32'h20c664b0
	         : (byte_in == 8'hd6)? 32'he0f5444e
	         : (byte_in == 8'hd7)? 32'h1c12624c
	         : (byte_in == 8'hd8)? 32'h5c46034f
	         : (byte_in == 8'hd9)? 32'ha0a1254d
	         : (byte_in == 8'hda)? 32'h609205b3
	         : (byte_in == 8'hdb)? 32'h9c7523b1
	         : (byte_in == 8'hdc)? 32'ha5884f4b
	         : (byte_in == 8'hdd)? 32'h596f6949
	         : (byte_in == 8'hde)? 32'h995c49b7
	         : (byte_in == 8'hdf)? 32'h65bb6fb5
	         : (byte_in == 8'he0)? 32'h4ed6c5e9
	         : (byte_in == 8'he1)? 32'hb231e3eb
	         : (byte_in == 8'he2)? 32'h7202c315
	         : (byte_in == 8'he3)? 32'h8ee5e517
	         : (byte_in == 8'he4)? 32'hb71889ed
	         : (byte_in == 8'he5)? 32'h4bffafef
	         : (byte_in == 8'he6)? 32'h8bcc8f11
	         : (byte_in == 8'he7)? 32'h772ba913
	         : (byte_in == 8'he8)? 32'h377fc810
	         : (byte_in == 8'he9)? 32'hcb98ee12
	         : (byte_in == 8'hea)? 32'h0babceec
	         : (byte_in == 8'heb)? 32'hf74ce8ee
	         : (byte_in == 8'hec)? 32'hceb18414
	         : (byte_in == 8'hed)? 32'h3256a216
	         : (byte_in == 8'hee)? 32'hf26582e8
	         : (byte_in == 8'hef)? 32'h0e82a4ea
	         : (byte_in == 8'hf0)? 32'h78b3ae41
	         : (byte_in == 8'hf1)? 32'h84548843
	         : (byte_in == 8'hf2)? 32'h4467a8bd
	         : (byte_in == 8'hf3)? 32'hb8808ebf
	         : (byte_in == 8'hf4)? 32'h817de245
	         : (byte_in == 8'hf5)? 32'h7d9ac447
	         : (byte_in == 8'hf6)? 32'hbda9e4b9
	         : (byte_in == 8'hf7)? 32'h414ec2bb
	         : (byte_in == 8'hf8)? 32'h011aa3b8
	         : (byte_in == 8'hf9)? 32'hfdfd85ba
	         : (byte_in == 8'hfa)? 32'h3dcea544
	         : (byte_in == 8'hfb)? 32'hc1298346
	         : (byte_in == 8'hfc)? 32'hf8d4efbc
	         : (byte_in == 8'hfd)? 32'h0433c9be
	         : (byte_in == 8'hfe)? 32'hc400e940
	         :                     32'h38e7cf42;

endmodule
//}}}

module TABLE10(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h8589d8ab
	         : (byte_in == 8'h02)? 32'ha29d1297
	         : (byte_in == 8'h03)? 32'h2714ca3c
	         : (byte_in == 8'h04)? 32'h60e5f9f2
	         : (byte_in == 8'h05)? 32'he56c2159
	         : (byte_in == 8'h06)? 32'hc278eb65
	         : (byte_in == 8'h07)? 32'h47f133ce
	         : (byte_in == 8'h08)? 32'h80c2d68f
	         : (byte_in == 8'h09)? 32'h054b0e24
	         : (byte_in == 8'h0a)? 32'h225fc418
	         : (byte_in == 8'h0b)? 32'ha7d61cb3
	         : (byte_in == 8'h0c)? 32'he0272f7d
	         : (byte_in == 8'h0d)? 32'h65aef7d6
	         : (byte_in == 8'h0e)? 32'h42ba3dea
	         : (byte_in == 8'h0f)? 32'hc733e541
	         : (byte_in == 8'h10)? 32'h6fc548e1
	         : (byte_in == 8'h11)? 32'hea4c904a
	         : (byte_in == 8'h12)? 32'hcd585a76
	         : (byte_in == 8'h13)? 32'h48d182dd
	         : (byte_in == 8'h14)? 32'h0f20b113
	         : (byte_in == 8'h15)? 32'h8aa969b8
	         : (byte_in == 8'h16)? 32'hadbda384
	         : (byte_in == 8'h17)? 32'h28347b2f
	         : (byte_in == 8'h18)? 32'hef079e6e
	         : (byte_in == 8'h19)? 32'h6a8e46c5
	         : (byte_in == 8'h1a)? 32'h4d9a8cf9
	         : (byte_in == 8'h1b)? 32'hc8135452
	         : (byte_in == 8'h1c)? 32'h8fe2679c
	         : (byte_in == 8'h1d)? 32'h0a6bbf37
	         : (byte_in == 8'h1e)? 32'h2d7f750b
	         : (byte_in == 8'h1f)? 32'ha8f6ada0
	         : (byte_in == 8'h20)? 32'h6a72e5bb
	         : (byte_in == 8'h21)? 32'heffb3d10
	         : (byte_in == 8'h22)? 32'hc8eff72c
	         : (byte_in == 8'h23)? 32'h4d662f87
	         : (byte_in == 8'h24)? 32'h0a971c49
	         : (byte_in == 8'h25)? 32'h8f1ec4e2
	         : (byte_in == 8'h26)? 32'ha80a0ede
	         : (byte_in == 8'h27)? 32'h2d83d675
	         : (byte_in == 8'h28)? 32'heab03334
	         : (byte_in == 8'h29)? 32'h6f39eb9f
	         : (byte_in == 8'h2a)? 32'h482d21a3
	         : (byte_in == 8'h2b)? 32'hcda4f908
	         : (byte_in == 8'h2c)? 32'h8a55cac6
	         : (byte_in == 8'h2d)? 32'h0fdc126d
	         : (byte_in == 8'h2e)? 32'h28c8d851
	         : (byte_in == 8'h2f)? 32'had4100fa
	         : (byte_in == 8'h30)? 32'h05b7ad5a
	         : (byte_in == 8'h31)? 32'h803e75f1
	         : (byte_in == 8'h32)? 32'ha72abfcd
	         : (byte_in == 8'h33)? 32'h22a36766
	         : (byte_in == 8'h34)? 32'h655254a8
	         : (byte_in == 8'h35)? 32'he0db8c03
	         : (byte_in == 8'h36)? 32'hc7cf463f
	         : (byte_in == 8'h37)? 32'h42469e94
	         : (byte_in == 8'h38)? 32'h85757bd5
	         : (byte_in == 8'h39)? 32'h00fca37e
	         : (byte_in == 8'h3a)? 32'h27e86942
	         : (byte_in == 8'h3b)? 32'ha261b1e9
	         : (byte_in == 8'h3c)? 32'he5908227
	         : (byte_in == 8'h3d)? 32'h60195a8c
	         : (byte_in == 8'h3e)? 32'h470d90b0
	         : (byte_in == 8'h3f)? 32'hc284481b
	         : (byte_in == 8'h40)? 32'h71852ac7
	         : (byte_in == 8'h41)? 32'hf40cf26c
	         : (byte_in == 8'h42)? 32'hd3183850
	         : (byte_in == 8'h43)? 32'h5691e0fb
	         : (byte_in == 8'h44)? 32'h1160d335
	         : (byte_in == 8'h45)? 32'h94e90b9e
	         : (byte_in == 8'h46)? 32'hb3fdc1a2
	         : (byte_in == 8'h47)? 32'h36741909
	         : (byte_in == 8'h48)? 32'hf147fc48
	         : (byte_in == 8'h49)? 32'h74ce24e3
	         : (byte_in == 8'h4a)? 32'h53daeedf
	         : (byte_in == 8'h4b)? 32'hd6533674
	         : (byte_in == 8'h4c)? 32'h91a205ba
	         : (byte_in == 8'h4d)? 32'h142bdd11
	         : (byte_in == 8'h4e)? 32'h333f172d
	         : (byte_in == 8'h4f)? 32'hb6b6cf86
	         : (byte_in == 8'h50)? 32'h1e406226
	         : (byte_in == 8'h51)? 32'h9bc9ba8d
	         : (byte_in == 8'h52)? 32'hbcdd70b1
	         : (byte_in == 8'h53)? 32'h3954a81a
	         : (byte_in == 8'h54)? 32'h7ea59bd4
	         : (byte_in == 8'h55)? 32'hfb2c437f
	         : (byte_in == 8'h56)? 32'hdc388943
	         : (byte_in == 8'h57)? 32'h59b151e8
	         : (byte_in == 8'h58)? 32'h9e82b4a9
	         : (byte_in == 8'h59)? 32'h1b0b6c02
	         : (byte_in == 8'h5a)? 32'h3c1fa63e
	         : (byte_in == 8'h5b)? 32'hb9967e95
	         : (byte_in == 8'h5c)? 32'hfe674d5b
	         : (byte_in == 8'h5d)? 32'h7bee95f0
	         : (byte_in == 8'h5e)? 32'h5cfa5fcc
	         : (byte_in == 8'h5f)? 32'hd9738767
	         : (byte_in == 8'h60)? 32'h1bf7cf7c
	         : (byte_in == 8'h61)? 32'h9e7e17d7
	         : (byte_in == 8'h62)? 32'hb96addeb
	         : (byte_in == 8'h63)? 32'h3ce30540
	         : (byte_in == 8'h64)? 32'h7b12368e
	         : (byte_in == 8'h65)? 32'hfe9bee25
	         : (byte_in == 8'h66)? 32'hd98f2419
	         : (byte_in == 8'h67)? 32'h5c06fcb2
	         : (byte_in == 8'h68)? 32'h9b3519f3
	         : (byte_in == 8'h69)? 32'h1ebcc158
	         : (byte_in == 8'h6a)? 32'h39a80b64
	         : (byte_in == 8'h6b)? 32'hbc21d3cf
	         : (byte_in == 8'h6c)? 32'hfbd0e001
	         : (byte_in == 8'h6d)? 32'h7e5938aa
	         : (byte_in == 8'h6e)? 32'h594df296
	         : (byte_in == 8'h6f)? 32'hdcc42a3d
	         : (byte_in == 8'h70)? 32'h7432879d
	         : (byte_in == 8'h71)? 32'hf1bb5f36
	         : (byte_in == 8'h72)? 32'hd6af950a
	         : (byte_in == 8'h73)? 32'h53264da1
	         : (byte_in == 8'h74)? 32'h14d77e6f
	         : (byte_in == 8'h75)? 32'h915ea6c4
	         : (byte_in == 8'h76)? 32'hb64a6cf8
	         : (byte_in == 8'h77)? 32'h33c3b453
	         : (byte_in == 8'h78)? 32'hf4f05112
	         : (byte_in == 8'h79)? 32'h717989b9
	         : (byte_in == 8'h7a)? 32'h566d4385
	         : (byte_in == 8'h7b)? 32'hd3e49b2e
	         : (byte_in == 8'h7c)? 32'h9415a8e0
	         : (byte_in == 8'h7d)? 32'h119c704b
	         : (byte_in == 8'h7e)? 32'h3688ba77
	         : (byte_in == 8'h7f)? 32'hb30162dc
	         : (byte_in == 8'h80)? 32'hbf1283d3
	         : (byte_in == 8'h81)? 32'h3a9b5b78
	         : (byte_in == 8'h82)? 32'h1d8f9144
	         : (byte_in == 8'h83)? 32'h980649ef
	         : (byte_in == 8'h84)? 32'hdff77a21
	         : (byte_in == 8'h85)? 32'h5a7ea28a
	         : (byte_in == 8'h86)? 32'h7d6a68b6
	         : (byte_in == 8'h87)? 32'hf8e3b01d
	         : (byte_in == 8'h88)? 32'h3fd0555c
	         : (byte_in == 8'h89)? 32'hba598df7
	         : (byte_in == 8'h8a)? 32'h9d4d47cb
	         : (byte_in == 8'h8b)? 32'h18c49f60
	         : (byte_in == 8'h8c)? 32'h5f35acae
	         : (byte_in == 8'h8d)? 32'hdabc7405
	         : (byte_in == 8'h8e)? 32'hfda8be39
	         : (byte_in == 8'h8f)? 32'h78216692
	         : (byte_in == 8'h90)? 32'hd0d7cb32
	         : (byte_in == 8'h91)? 32'h555e1399
	         : (byte_in == 8'h92)? 32'h724ad9a5
	         : (byte_in == 8'h93)? 32'hf7c3010e
	         : (byte_in == 8'h94)? 32'hb03232c0
	         : (byte_in == 8'h95)? 32'h35bbea6b
	         : (byte_in == 8'h96)? 32'h12af2057
	         : (byte_in == 8'h97)? 32'h9726f8fc
	         : (byte_in == 8'h98)? 32'h50151dbd
	         : (byte_in == 8'h99)? 32'hd59cc516
	         : (byte_in == 8'h9a)? 32'hf2880f2a
	         : (byte_in == 8'h9b)? 32'h7701d781
	         : (byte_in == 8'h9c)? 32'h30f0e44f
	         : (byte_in == 8'h9d)? 32'hb5793ce4
	         : (byte_in == 8'h9e)? 32'h926df6d8
	         : (byte_in == 8'h9f)? 32'h17e42e73
	         : (byte_in == 8'ha0)? 32'hd5606668
	         : (byte_in == 8'ha1)? 32'h50e9bec3
	         : (byte_in == 8'ha2)? 32'h77fd74ff
	         : (byte_in == 8'ha3)? 32'hf274ac54
	         : (byte_in == 8'ha4)? 32'hb5859f9a
	         : (byte_in == 8'ha5)? 32'h300c4731
	         : (byte_in == 8'ha6)? 32'h17188d0d
	         : (byte_in == 8'ha7)? 32'h929155a6
	         : (byte_in == 8'ha8)? 32'h55a2b0e7
	         : (byte_in == 8'ha9)? 32'hd02b684c
	         : (byte_in == 8'haa)? 32'hf73fa270
	         : (byte_in == 8'hab)? 32'h72b67adb
	         : (byte_in == 8'hac)? 32'h35474915
	         : (byte_in == 8'had)? 32'hb0ce91be
	         : (byte_in == 8'hae)? 32'h97da5b82
	         : (byte_in == 8'haf)? 32'h12538329
	         : (byte_in == 8'hb0)? 32'hbaa52e89
	         : (byte_in == 8'hb1)? 32'h3f2cf622
	         : (byte_in == 8'hb2)? 32'h18383c1e
	         : (byte_in == 8'hb3)? 32'h9db1e4b5
	         : (byte_in == 8'hb4)? 32'hda40d77b
	         : (byte_in == 8'hb5)? 32'h5fc90fd0
	         : (byte_in == 8'hb6)? 32'h78ddc5ec
	         : (byte_in == 8'hb7)? 32'hfd541d47
	         : (byte_in == 8'hb8)? 32'h3a67f806
	         : (byte_in == 8'hb9)? 32'hbfee20ad
	         : (byte_in == 8'hba)? 32'h98faea91
	         : (byte_in == 8'hbb)? 32'h1d73323a
	         : (byte_in == 8'hbc)? 32'h5a8201f4
	         : (byte_in == 8'hbd)? 32'hdf0bd95f
	         : (byte_in == 8'hbe)? 32'hf81f1363
	         : (byte_in == 8'hbf)? 32'h7d96cbc8
	         : (byte_in == 8'hc0)? 32'hce97a914
	         : (byte_in == 8'hc1)? 32'h4b1e71bf
	         : (byte_in == 8'hc2)? 32'h6c0abb83
	         : (byte_in == 8'hc3)? 32'he9836328
	         : (byte_in == 8'hc4)? 32'hae7250e6
	         : (byte_in == 8'hc5)? 32'h2bfb884d
	         : (byte_in == 8'hc6)? 32'h0cef4271
	         : (byte_in == 8'hc7)? 32'h89669ada
	         : (byte_in == 8'hc8)? 32'h4e557f9b
	         : (byte_in == 8'hc9)? 32'hcbdca730
	         : (byte_in == 8'hca)? 32'hecc86d0c
	         : (byte_in == 8'hcb)? 32'h6941b5a7
	         : (byte_in == 8'hcc)? 32'h2eb08669
	         : (byte_in == 8'hcd)? 32'hab395ec2
	         : (byte_in == 8'hce)? 32'h8c2d94fe
	         : (byte_in == 8'hcf)? 32'h09a44c55
	         : (byte_in == 8'hd0)? 32'ha152e1f5
	         : (byte_in == 8'hd1)? 32'h24db395e
	         : (byte_in == 8'hd2)? 32'h03cff362
	         : (byte_in == 8'hd3)? 32'h86462bc9
	         : (byte_in == 8'hd4)? 32'hc1b71807
	         : (byte_in == 8'hd5)? 32'h443ec0ac
	         : (byte_in == 8'hd6)? 32'h632a0a90
	         : (byte_in == 8'hd7)? 32'he6a3d23b
	         : (byte_in == 8'hd8)? 32'h2190377a
	         : (byte_in == 8'hd9)? 32'ha419efd1
	         : (byte_in == 8'hda)? 32'h830d25ed
	         : (byte_in == 8'hdb)? 32'h0684fd46
	         : (byte_in == 8'hdc)? 32'h4175ce88
	         : (byte_in == 8'hdd)? 32'hc4fc1623
	         : (byte_in == 8'hde)? 32'he3e8dc1f
	         : (byte_in == 8'hdf)? 32'h666104b4
	         : (byte_in == 8'he0)? 32'ha4e54caf
	         : (byte_in == 8'he1)? 32'h216c9404
	         : (byte_in == 8'he2)? 32'h06785e38
	         : (byte_in == 8'he3)? 32'h83f18693
	         : (byte_in == 8'he4)? 32'hc400b55d
	         : (byte_in == 8'he5)? 32'h41896df6
	         : (byte_in == 8'he6)? 32'h669da7ca
	         : (byte_in == 8'he7)? 32'he3147f61
	         : (byte_in == 8'he8)? 32'h24279a20
	         : (byte_in == 8'he9)? 32'ha1ae428b
	         : (byte_in == 8'hea)? 32'h86ba88b7
	         : (byte_in == 8'heb)? 32'h0333501c
	         : (byte_in == 8'hec)? 32'h44c263d2
	         : (byte_in == 8'hed)? 32'hc14bbb79
	         : (byte_in == 8'hee)? 32'he65f7145
	         : (byte_in == 8'hef)? 32'h63d6a9ee
	         : (byte_in == 8'hf0)? 32'hcb20044e
	         : (byte_in == 8'hf1)? 32'h4ea9dce5
	         : (byte_in == 8'hf2)? 32'h69bd16d9
	         : (byte_in == 8'hf3)? 32'hec34ce72
	         : (byte_in == 8'hf4)? 32'habc5fdbc
	         : (byte_in == 8'hf5)? 32'h2e4c2517
	         : (byte_in == 8'hf6)? 32'h0958ef2b
	         : (byte_in == 8'hf7)? 32'h8cd13780
	         : (byte_in == 8'hf8)? 32'h4be2d2c1
	         : (byte_in == 8'hf9)? 32'hce6b0a6a
	         : (byte_in == 8'hfa)? 32'he97fc056
	         : (byte_in == 8'hfb)? 32'h6cf618fd
	         : (byte_in == 8'hfc)? 32'h2b072b33
	         : (byte_in == 8'hfd)? 32'hae8ef398
	         : (byte_in == 8'hfe)? 32'h899a39a4
	         :                     32'h0c13e10f;

endmodule
//}}}

module TABLE11(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h88fd1d2b
	         : (byte_in == 8'h02)? 32'hbbdcf407
	         : (byte_in == 8'h03)? 32'h3321e92c
	         : (byte_in == 8'h04)? 32'h11fa3a57
	         : (byte_in == 8'h05)? 32'h9907277c
	         : (byte_in == 8'h06)? 32'haa26ce50
	         : (byte_in == 8'h07)? 32'h22dbd37b
	         : (byte_in == 8'h08)? 32'h77b9e80f
	         : (byte_in == 8'h09)? 32'hff44f524
	         : (byte_in == 8'h0a)? 32'hcc651c08
	         : (byte_in == 8'h0b)? 32'h44980123
	         : (byte_in == 8'h0c)? 32'h6643d258
	         : (byte_in == 8'h0d)? 32'heebecf73
	         : (byte_in == 8'h0e)? 32'hdd9f265f
	         : (byte_in == 8'h0f)? 32'h55623b74
	         : (byte_in == 8'h10)? 32'h8dfacfab
	         : (byte_in == 8'h11)? 32'h0507d280
	         : (byte_in == 8'h12)? 32'h36263bac
	         : (byte_in == 8'h13)? 32'hbedb2687
	         : (byte_in == 8'h14)? 32'h9c00f5fc
	         : (byte_in == 8'h15)? 32'h14fde8d7
	         : (byte_in == 8'h16)? 32'h27dc01fb
	         : (byte_in == 8'h17)? 32'haf211cd0
	         : (byte_in == 8'h18)? 32'hfa4327a4
	         : (byte_in == 8'h19)? 32'h72be3a8f
	         : (byte_in == 8'h1a)? 32'h419fd3a3
	         : (byte_in == 8'h1b)? 32'hc962ce88
	         : (byte_in == 8'h1c)? 32'hebb91df3
	         : (byte_in == 8'h1d)? 32'h634400d8
	         : (byte_in == 8'h1e)? 32'h5065e9f4
	         : (byte_in == 8'h1f)? 32'hd898f4df
	         : (byte_in == 8'h20)? 32'h848598ba
	         : (byte_in == 8'h21)? 32'h0c788591
	         : (byte_in == 8'h22)? 32'h3f596cbd
	         : (byte_in == 8'h23)? 32'hb7a47196
	         : (byte_in == 8'h24)? 32'h957fa2ed
	         : (byte_in == 8'h25)? 32'h1d82bfc6
	         : (byte_in == 8'h26)? 32'h2ea356ea
	         : (byte_in == 8'h27)? 32'ha65e4bc1
	         : (byte_in == 8'h28)? 32'hf33c70b5
	         : (byte_in == 8'h29)? 32'h7bc16d9e
	         : (byte_in == 8'h2a)? 32'h48e084b2
	         : (byte_in == 8'h2b)? 32'hc01d9999
	         : (byte_in == 8'h2c)? 32'he2c64ae2
	         : (byte_in == 8'h2d)? 32'h6a3b57c9
	         : (byte_in == 8'h2e)? 32'h591abee5
	         : (byte_in == 8'h2f)? 32'hd1e7a3ce
	         : (byte_in == 8'h30)? 32'h097f5711
	         : (byte_in == 8'h31)? 32'h81824a3a
	         : (byte_in == 8'h32)? 32'hb2a3a316
	         : (byte_in == 8'h33)? 32'h3a5ebe3d
	         : (byte_in == 8'h34)? 32'h18856d46
	         : (byte_in == 8'h35)? 32'h9078706d
	         : (byte_in == 8'h36)? 32'ha3599941
	         : (byte_in == 8'h37)? 32'h2ba4846a
	         : (byte_in == 8'h38)? 32'h7ec6bf1e
	         : (byte_in == 8'h39)? 32'hf63ba235
	         : (byte_in == 8'h3a)? 32'hc51a4b19
	         : (byte_in == 8'h3b)? 32'h4de75632
	         : (byte_in == 8'h3c)? 32'h6f3c8549
	         : (byte_in == 8'h3d)? 32'he7c19862
	         : (byte_in == 8'h3e)? 32'hd4e0714e
	         : (byte_in == 8'h3f)? 32'h5c1d6c65
	         : (byte_in == 8'h40)? 32'hb5fb2452
	         : (byte_in == 8'h41)? 32'h3d063979
	         : (byte_in == 8'h42)? 32'h0e27d055
	         : (byte_in == 8'h43)? 32'h86dacd7e
	         : (byte_in == 8'h44)? 32'ha4011e05
	         : (byte_in == 8'h45)? 32'h2cfc032e
	         : (byte_in == 8'h46)? 32'h1fddea02
	         : (byte_in == 8'h47)? 32'h9720f729
	         : (byte_in == 8'h48)? 32'hc242cc5d
	         : (byte_in == 8'h49)? 32'h4abfd176
	         : (byte_in == 8'h4a)? 32'h799e385a
	         : (byte_in == 8'h4b)? 32'hf1632571
	         : (byte_in == 8'h4c)? 32'hd3b8f60a
	         : (byte_in == 8'h4d)? 32'h5b45eb21
	         : (byte_in == 8'h4e)? 32'h6864020d
	         : (byte_in == 8'h4f)? 32'he0991f26
	         : (byte_in == 8'h50)? 32'h3801ebf9
	         : (byte_in == 8'h51)? 32'hb0fcf6d2
	         : (byte_in == 8'h52)? 32'h83dd1ffe
	         : (byte_in == 8'h53)? 32'h0b2002d5
	         : (byte_in == 8'h54)? 32'h29fbd1ae
	         : (byte_in == 8'h55)? 32'ha106cc85
	         : (byte_in == 8'h56)? 32'h922725a9
	         : (byte_in == 8'h57)? 32'h1ada3882
	         : (byte_in == 8'h58)? 32'h4fb803f6
	         : (byte_in == 8'h59)? 32'hc7451edd
	         : (byte_in == 8'h5a)? 32'hf464f7f1
	         : (byte_in == 8'h5b)? 32'h7c99eada
	         : (byte_in == 8'h5c)? 32'h5e4239a1
	         : (byte_in == 8'h5d)? 32'hd6bf248a
	         : (byte_in == 8'h5e)? 32'he59ecda6
	         : (byte_in == 8'h5f)? 32'h6d63d08d
	         : (byte_in == 8'h60)? 32'h317ebce8
	         : (byte_in == 8'h61)? 32'hb983a1c3
	         : (byte_in == 8'h62)? 32'h8aa248ef
	         : (byte_in == 8'h63)? 32'h025f55c4
	         : (byte_in == 8'h64)? 32'h208486bf
	         : (byte_in == 8'h65)? 32'ha8799b94
	         : (byte_in == 8'h66)? 32'h9b5872b8
	         : (byte_in == 8'h67)? 32'h13a56f93
	         : (byte_in == 8'h68)? 32'h46c754e7
	         : (byte_in == 8'h69)? 32'hce3a49cc
	         : (byte_in == 8'h6a)? 32'hfd1ba0e0
	         : (byte_in == 8'h6b)? 32'h75e6bdcb
	         : (byte_in == 8'h6c)? 32'h573d6eb0
	         : (byte_in == 8'h6d)? 32'hdfc0739b
	         : (byte_in == 8'h6e)? 32'hece19ab7
	         : (byte_in == 8'h6f)? 32'h641c879c
	         : (byte_in == 8'h70)? 32'hbc847343
	         : (byte_in == 8'h71)? 32'h34796e68
	         : (byte_in == 8'h72)? 32'h07588744
	         : (byte_in == 8'h73)? 32'h8fa59a6f
	         : (byte_in == 8'h74)? 32'had7e4914
	         : (byte_in == 8'h75)? 32'h2583543f
	         : (byte_in == 8'h76)? 32'h16a2bd13
	         : (byte_in == 8'h77)? 32'h9e5fa038
	         : (byte_in == 8'h78)? 32'hcb3d9b4c
	         : (byte_in == 8'h79)? 32'h43c08667
	         : (byte_in == 8'h7a)? 32'h70e16f4b
	         : (byte_in == 8'h7b)? 32'hf81c7260
	         : (byte_in == 8'h7c)? 32'hdac7a11b
	         : (byte_in == 8'h7d)? 32'h523abc30
	         : (byte_in == 8'h7e)? 32'h611b551c
	         : (byte_in == 8'h7f)? 32'he9e64837
	         : (byte_in == 8'h80)? 32'h62fc79d0
	         : (byte_in == 8'h81)? 32'hea0164fb
	         : (byte_in == 8'h82)? 32'hd9208dd7
	         : (byte_in == 8'h83)? 32'h51dd90fc
	         : (byte_in == 8'h84)? 32'h73064387
	         : (byte_in == 8'h85)? 32'hfbfb5eac
	         : (byte_in == 8'h86)? 32'hc8dab780
	         : (byte_in == 8'h87)? 32'h4027aaab
	         : (byte_in == 8'h88)? 32'h154591df
	         : (byte_in == 8'h89)? 32'h9db88cf4
	         : (byte_in == 8'h8a)? 32'hae9965d8
	         : (byte_in == 8'h8b)? 32'h266478f3
	         : (byte_in == 8'h8c)? 32'h04bfab88
	         : (byte_in == 8'h8d)? 32'h8c42b6a3
	         : (byte_in == 8'h8e)? 32'hbf635f8f
	         : (byte_in == 8'h8f)? 32'h379e42a4
	         : (byte_in == 8'h90)? 32'hef06b67b
	         : (byte_in == 8'h91)? 32'h67fbab50
	         : (byte_in == 8'h92)? 32'h54da427c
	         : (byte_in == 8'h93)? 32'hdc275f57
	         : (byte_in == 8'h94)? 32'hfefc8c2c
	         : (byte_in == 8'h95)? 32'h76019107
	         : (byte_in == 8'h96)? 32'h4520782b
	         : (byte_in == 8'h97)? 32'hcddd6500
	         : (byte_in == 8'h98)? 32'h98bf5e74
	         : (byte_in == 8'h99)? 32'h1042435f
	         : (byte_in == 8'h9a)? 32'h2363aa73
	         : (byte_in == 8'h9b)? 32'hab9eb758
	         : (byte_in == 8'h9c)? 32'h89456423
	         : (byte_in == 8'h9d)? 32'h01b87908
	         : (byte_in == 8'h9e)? 32'h32999024
	         : (byte_in == 8'h9f)? 32'hba648d0f
	         : (byte_in == 8'ha0)? 32'he679e16a
	         : (byte_in == 8'ha1)? 32'h6e84fc41
	         : (byte_in == 8'ha2)? 32'h5da5156d
	         : (byte_in == 8'ha3)? 32'hd5580846
	         : (byte_in == 8'ha4)? 32'hf783db3d
	         : (byte_in == 8'ha5)? 32'h7f7ec616
	         : (byte_in == 8'ha6)? 32'h4c5f2f3a
	         : (byte_in == 8'ha7)? 32'hc4a23211
	         : (byte_in == 8'ha8)? 32'h91c00965
	         : (byte_in == 8'ha9)? 32'h193d144e
	         : (byte_in == 8'haa)? 32'h2a1cfd62
	         : (byte_in == 8'hab)? 32'ha2e1e049
	         : (byte_in == 8'hac)? 32'h803a3332
	         : (byte_in == 8'had)? 32'h08c72e19
	         : (byte_in == 8'hae)? 32'h3be6c735
	         : (byte_in == 8'haf)? 32'hb31bda1e
	         : (byte_in == 8'hb0)? 32'h6b832ec1
	         : (byte_in == 8'hb1)? 32'he37e33ea
	         : (byte_in == 8'hb2)? 32'hd05fdac6
	         : (byte_in == 8'hb3)? 32'h58a2c7ed
	         : (byte_in == 8'hb4)? 32'h7a791496
	         : (byte_in == 8'hb5)? 32'hf28409bd
	         : (byte_in == 8'hb6)? 32'hc1a5e091
	         : (byte_in == 8'hb7)? 32'h4958fdba
	         : (byte_in == 8'hb8)? 32'h1c3ac6ce
	         : (byte_in == 8'hb9)? 32'h94c7dbe5
	         : (byte_in == 8'hba)? 32'ha7e632c9
	         : (byte_in == 8'hbb)? 32'h2f1b2fe2
	         : (byte_in == 8'hbc)? 32'h0dc0fc99
	         : (byte_in == 8'hbd)? 32'h853de1b2
	         : (byte_in == 8'hbe)? 32'hb61c089e
	         : (byte_in == 8'hbf)? 32'h3ee115b5
	         : (byte_in == 8'hc0)? 32'hd7075d82
	         : (byte_in == 8'hc1)? 32'h5ffa40a9
	         : (byte_in == 8'hc2)? 32'h6cdba985
	         : (byte_in == 8'hc3)? 32'he426b4ae
	         : (byte_in == 8'hc4)? 32'hc6fd67d5
	         : (byte_in == 8'hc5)? 32'h4e007afe
	         : (byte_in == 8'hc6)? 32'h7d2193d2
	         : (byte_in == 8'hc7)? 32'hf5dc8ef9
	         : (byte_in == 8'hc8)? 32'ha0beb58d
	         : (byte_in == 8'hc9)? 32'h2843a8a6
	         : (byte_in == 8'hca)? 32'h1b62418a
	         : (byte_in == 8'hcb)? 32'h939f5ca1
	         : (byte_in == 8'hcc)? 32'hb1448fda
	         : (byte_in == 8'hcd)? 32'h39b992f1
	         : (byte_in == 8'hce)? 32'h0a987bdd
	         : (byte_in == 8'hcf)? 32'h826566f6
	         : (byte_in == 8'hd0)? 32'h5afd9229
	         : (byte_in == 8'hd1)? 32'hd2008f02
	         : (byte_in == 8'hd2)? 32'he121662e
	         : (byte_in == 8'hd3)? 32'h69dc7b05
	         : (byte_in == 8'hd4)? 32'h4b07a87e
	         : (byte_in == 8'hd5)? 32'hc3fab555
	         : (byte_in == 8'hd6)? 32'hf0db5c79
	         : (byte_in == 8'hd7)? 32'h78264152
	         : (byte_in == 8'hd8)? 32'h2d447a26
	         : (byte_in == 8'hd9)? 32'ha5b9670d
	         : (byte_in == 8'hda)? 32'h96988e21
	         : (byte_in == 8'hdb)? 32'h1e65930a
	         : (byte_in == 8'hdc)? 32'h3cbe4071
	         : (byte_in == 8'hdd)? 32'hb4435d5a
	         : (byte_in == 8'hde)? 32'h8762b476
	         : (byte_in == 8'hdf)? 32'h0f9fa95d
	         : (byte_in == 8'he0)? 32'h5382c538
	         : (byte_in == 8'he1)? 32'hdb7fd813
	         : (byte_in == 8'he2)? 32'he85e313f
	         : (byte_in == 8'he3)? 32'h60a32c14
	         : (byte_in == 8'he4)? 32'h4278ff6f
	         : (byte_in == 8'he5)? 32'hca85e244
	         : (byte_in == 8'he6)? 32'hf9a40b68
	         : (byte_in == 8'he7)? 32'h71591643
	         : (byte_in == 8'he8)? 32'h243b2d37
	         : (byte_in == 8'he9)? 32'hacc6301c
	         : (byte_in == 8'hea)? 32'h9fe7d930
	         : (byte_in == 8'heb)? 32'h171ac41b
	         : (byte_in == 8'hec)? 32'h35c11760
	         : (byte_in == 8'hed)? 32'hbd3c0a4b
	         : (byte_in == 8'hee)? 32'h8e1de367
	         : (byte_in == 8'hef)? 32'h06e0fe4c
	         : (byte_in == 8'hf0)? 32'hde780a93
	         : (byte_in == 8'hf1)? 32'h568517b8
	         : (byte_in == 8'hf2)? 32'h65a4fe94
	         : (byte_in == 8'hf3)? 32'hed59e3bf
	         : (byte_in == 8'hf4)? 32'hcf8230c4
	         : (byte_in == 8'hf5)? 32'h477f2def
	         : (byte_in == 8'hf6)? 32'h745ec4c3
	         : (byte_in == 8'hf7)? 32'hfca3d9e8
	         : (byte_in == 8'hf8)? 32'ha9c1e29c
	         : (byte_in == 8'hf9)? 32'h213cffb7
	         : (byte_in == 8'hfa)? 32'h121d169b
	         : (byte_in == 8'hfb)? 32'h9ae00bb0
	         : (byte_in == 8'hfc)? 32'hb83bd8cb
	         : (byte_in == 8'hfd)? 32'h30c6c5e0
	         : (byte_in == 8'hfe)? 32'h03e72ccc
	         :                     32'h8b1a31e7;

endmodule
//}}}

module TABLE12(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'hb5a4c63b
	         : (byte_in == 8'h02)? 32'h539cbdbf
	         : (byte_in == 8'h03)? 32'he6387b84
	         : (byte_in == 8'h04)? 32'h8d75f7f1
	         : (byte_in == 8'h05)? 32'h38d131ca
	         : (byte_in == 8'h06)? 32'hdee94a4e
	         : (byte_in == 8'h07)? 32'h6b4d8c75
	         : (byte_in == 8'h08)? 32'h1298bd46
	         : (byte_in == 8'h09)? 32'ha73c7b7d
	         : (byte_in == 8'h0a)? 32'h410400f9
	         : (byte_in == 8'h0b)? 32'hf4a0c6c2
	         : (byte_in == 8'h0c)? 32'h9fed4ab7
	         : (byte_in == 8'h0d)? 32'h2a498c8c
	         : (byte_in == 8'h0e)? 32'hcc71f708
	         : (byte_in == 8'h0f)? 32'h79d53133
	         : (byte_in == 8'h10)? 32'haf4a29da
	         : (byte_in == 8'h11)? 32'h1aeeefe1
	         : (byte_in == 8'h12)? 32'hfcd69465
	         : (byte_in == 8'h13)? 32'h4972525e
	         : (byte_in == 8'h14)? 32'h223fde2b
	         : (byte_in == 8'h15)? 32'h979b1810
	         : (byte_in == 8'h16)? 32'h71a36394
	         : (byte_in == 8'h17)? 32'hc407a5af
	         : (byte_in == 8'h18)? 32'hbdd2949c
	         : (byte_in == 8'h19)? 32'h087652a7
	         : (byte_in == 8'h1a)? 32'hee4e2923
	         : (byte_in == 8'h1b)? 32'h5beaef18
	         : (byte_in == 8'h1c)? 32'h30a7636d
	         : (byte_in == 8'h1d)? 32'h8503a556
	         : (byte_in == 8'h1e)? 32'h633bded2
	         : (byte_in == 8'h1f)? 32'hd69f18e9
	         : (byte_in == 8'h20)? 32'h76acc733
	         : (byte_in == 8'h21)? 32'hc3080108
	         : (byte_in == 8'h22)? 32'h25307a8c
	         : (byte_in == 8'h23)? 32'h9094bcb7
	         : (byte_in == 8'h24)? 32'hfbd930c2
	         : (byte_in == 8'h25)? 32'h4e7df6f9
	         : (byte_in == 8'h26)? 32'ha8458d7d
	         : (byte_in == 8'h27)? 32'h1de14b46
	         : (byte_in == 8'h28)? 32'h64347a75
	         : (byte_in == 8'h29)? 32'hd190bc4e
	         : (byte_in == 8'h2a)? 32'h37a8c7ca
	         : (byte_in == 8'h2b)? 32'h820c01f1
	         : (byte_in == 8'h2c)? 32'he9418d84
	         : (byte_in == 8'h2d)? 32'h5ce54bbf
	         : (byte_in == 8'h2e)? 32'hbadd303b
	         : (byte_in == 8'h2f)? 32'h0f79f600
	         : (byte_in == 8'h30)? 32'hd9e6eee9
	         : (byte_in == 8'h31)? 32'h6c4228d2
	         : (byte_in == 8'h32)? 32'h8a7a5356
	         : (byte_in == 8'h33)? 32'h3fde956d
	         : (byte_in == 8'h34)? 32'h54931918
	         : (byte_in == 8'h35)? 32'he137df23
	         : (byte_in == 8'h36)? 32'h070fa4a7
	         : (byte_in == 8'h37)? 32'hb2ab629c
	         : (byte_in == 8'h38)? 32'hcb7e53af
	         : (byte_in == 8'h39)? 32'h7eda9594
	         : (byte_in == 8'h3a)? 32'h98e2ee10
	         : (byte_in == 8'h3b)? 32'h2d46282b
	         : (byte_in == 8'h3c)? 32'h460ba45e
	         : (byte_in == 8'h3d)? 32'hf3af6265
	         : (byte_in == 8'h3e)? 32'h159719e1
	         : (byte_in == 8'h3f)? 32'ha033dfda
	         : (byte_in == 8'h40)? 32'hb8a92831
	         : (byte_in == 8'h41)? 32'h0d0dee0a
	         : (byte_in == 8'h42)? 32'heb35958e
	         : (byte_in == 8'h43)? 32'h5e9153b5
	         : (byte_in == 8'h44)? 32'h35dcdfc0
	         : (byte_in == 8'h45)? 32'h807819fb
	         : (byte_in == 8'h46)? 32'h6640627f
	         : (byte_in == 8'h47)? 32'hd3e4a444
	         : (byte_in == 8'h48)? 32'haa319577
	         : (byte_in == 8'h49)? 32'h1f95534c
	         : (byte_in == 8'h4a)? 32'hf9ad28c8
	         : (byte_in == 8'h4b)? 32'h4c09eef3
	         : (byte_in == 8'h4c)? 32'h27446286
	         : (byte_in == 8'h4d)? 32'h92e0a4bd
	         : (byte_in == 8'h4e)? 32'h74d8df39
	         : (byte_in == 8'h4f)? 32'hc17c1902
	         : (byte_in == 8'h50)? 32'h17e301eb
	         : (byte_in == 8'h51)? 32'ha247c7d0
	         : (byte_in == 8'h52)? 32'h447fbc54
	         : (byte_in == 8'h53)? 32'hf1db7a6f
	         : (byte_in == 8'h54)? 32'h9a96f61a
	         : (byte_in == 8'h55)? 32'h2f323021
	         : (byte_in == 8'h56)? 32'hc90a4ba5
	         : (byte_in == 8'h57)? 32'h7cae8d9e
	         : (byte_in == 8'h58)? 32'h057bbcad
	         : (byte_in == 8'h59)? 32'hb0df7a96
	         : (byte_in == 8'h5a)? 32'h56e70112
	         : (byte_in == 8'h5b)? 32'he343c729
	         : (byte_in == 8'h5c)? 32'h880e4b5c
	         : (byte_in == 8'h5d)? 32'h3daa8d67
	         : (byte_in == 8'h5e)? 32'hdb92f6e3
	         : (byte_in == 8'h5f)? 32'h6e3630d8
	         : (byte_in == 8'h60)? 32'hce05ef02
	         : (byte_in == 8'h61)? 32'h7ba12939
	         : (byte_in == 8'h62)? 32'h9d9952bd
	         : (byte_in == 8'h63)? 32'h283d9486
	         : (byte_in == 8'h64)? 32'h437018f3
	         : (byte_in == 8'h65)? 32'hf6d4dec8
	         : (byte_in == 8'h66)? 32'h10eca54c
	         : (byte_in == 8'h67)? 32'ha5486377
	         : (byte_in == 8'h68)? 32'hdc9d5244
	         : (byte_in == 8'h69)? 32'h6939947f
	         : (byte_in == 8'h6a)? 32'h8f01effb
	         : (byte_in == 8'h6b)? 32'h3aa529c0
	         : (byte_in == 8'h6c)? 32'h51e8a5b5
	         : (byte_in == 8'h6d)? 32'he44c638e
	         : (byte_in == 8'h6e)? 32'h0274180a
	         : (byte_in == 8'h6f)? 32'hb7d0de31
	         : (byte_in == 8'h70)? 32'h614fc6d8
	         : (byte_in == 8'h71)? 32'hd4eb00e3
	         : (byte_in == 8'h72)? 32'h32d37b67
	         : (byte_in == 8'h73)? 32'h8777bd5c
	         : (byte_in == 8'h74)? 32'hec3a3129
	         : (byte_in == 8'h75)? 32'h599ef712
	         : (byte_in == 8'h76)? 32'hbfa68c96
	         : (byte_in == 8'h77)? 32'h0a024aad
	         : (byte_in == 8'h78)? 32'h73d77b9e
	         : (byte_in == 8'h79)? 32'hc673bda5
	         : (byte_in == 8'h7a)? 32'h204bc621
	         : (byte_in == 8'h7b)? 32'h95ef001a
	         : (byte_in == 8'h7c)? 32'hfea28c6f
	         : (byte_in == 8'h7d)? 32'h4b064a54
	         : (byte_in == 8'h7e)? 32'had3e31d0
	         : (byte_in == 8'h7f)? 32'h189af7eb
	         : (byte_in == 8'h80)? 32'h58f8485f
	         : (byte_in == 8'h81)? 32'hed5c8e64
	         : (byte_in == 8'h82)? 32'h0b64f5e0
	         : (byte_in == 8'h83)? 32'hbec033db
	         : (byte_in == 8'h84)? 32'hd58dbfae
	         : (byte_in == 8'h85)? 32'h60297995
	         : (byte_in == 8'h86)? 32'h86110211
	         : (byte_in == 8'h87)? 32'h33b5c42a
	         : (byte_in == 8'h88)? 32'h4a60f519
	         : (byte_in == 8'h89)? 32'hffc43322
	         : (byte_in == 8'h8a)? 32'h19fc48a6
	         : (byte_in == 8'h8b)? 32'hac588e9d
	         : (byte_in == 8'h8c)? 32'hc71502e8
	         : (byte_in == 8'h8d)? 32'h72b1c4d3
	         : (byte_in == 8'h8e)? 32'h9489bf57
	         : (byte_in == 8'h8f)? 32'h212d796c
	         : (byte_in == 8'h90)? 32'hf7b26185
	         : (byte_in == 8'h91)? 32'h4216a7be
	         : (byte_in == 8'h92)? 32'ha42edc3a
	         : (byte_in == 8'h93)? 32'h118a1a01
	         : (byte_in == 8'h94)? 32'h7ac79674
	         : (byte_in == 8'h95)? 32'hcf63504f
	         : (byte_in == 8'h96)? 32'h295b2bcb
	         : (byte_in == 8'h97)? 32'h9cffedf0
	         : (byte_in == 8'h98)? 32'he52adcc3
	         : (byte_in == 8'h99)? 32'h508e1af8
	         : (byte_in == 8'h9a)? 32'hb6b6617c
	         : (byte_in == 8'h9b)? 32'h0312a747
	         : (byte_in == 8'h9c)? 32'h685f2b32
	         : (byte_in == 8'h9d)? 32'hddfbed09
	         : (byte_in == 8'h9e)? 32'h3bc3968d
	         : (byte_in == 8'h9f)? 32'h8e6750b6
	         : (byte_in == 8'ha0)? 32'h2e548f6c
	         : (byte_in == 8'ha1)? 32'h9bf04957
	         : (byte_in == 8'ha2)? 32'h7dc832d3
	         : (byte_in == 8'ha3)? 32'hc86cf4e8
	         : (byte_in == 8'ha4)? 32'ha321789d
	         : (byte_in == 8'ha5)? 32'h1685bea6
	         : (byte_in == 8'ha6)? 32'hf0bdc522
	         : (byte_in == 8'ha7)? 32'h45190319
	         : (byte_in == 8'ha8)? 32'h3ccc322a
	         : (byte_in == 8'ha9)? 32'h8968f411
	         : (byte_in == 8'haa)? 32'h6f508f95
	         : (byte_in == 8'hab)? 32'hdaf449ae
	         : (byte_in == 8'hac)? 32'hb1b9c5db
	         : (byte_in == 8'had)? 32'h041d03e0
	         : (byte_in == 8'hae)? 32'he2257864
	         : (byte_in == 8'haf)? 32'h5781be5f
	         : (byte_in == 8'hb0)? 32'h811ea6b6
	         : (byte_in == 8'hb1)? 32'h34ba608d
	         : (byte_in == 8'hb2)? 32'hd2821b09
	         : (byte_in == 8'hb3)? 32'h6726dd32
	         : (byte_in == 8'hb4)? 32'h0c6b5147
	         : (byte_in == 8'hb5)? 32'hb9cf977c
	         : (byte_in == 8'hb6)? 32'h5ff7ecf8
	         : (byte_in == 8'hb7)? 32'hea532ac3
	         : (byte_in == 8'hb8)? 32'h93861bf0
	         : (byte_in == 8'hb9)? 32'h2622ddcb
	         : (byte_in == 8'hba)? 32'hc01aa64f
	         : (byte_in == 8'hbb)? 32'h75be6074
	         : (byte_in == 8'hbc)? 32'h1ef3ec01
	         : (byte_in == 8'hbd)? 32'hab572a3a
	         : (byte_in == 8'hbe)? 32'h4d6f51be
	         : (byte_in == 8'hbf)? 32'hf8cb9785
	         : (byte_in == 8'hc0)? 32'he051606e
	         : (byte_in == 8'hc1)? 32'h55f5a655
	         : (byte_in == 8'hc2)? 32'hb3cdddd1
	         : (byte_in == 8'hc3)? 32'h06691bea
	         : (byte_in == 8'hc4)? 32'h6d24979f
	         : (byte_in == 8'hc5)? 32'hd88051a4
	         : (byte_in == 8'hc6)? 32'h3eb82a20
	         : (byte_in == 8'hc7)? 32'h8b1cec1b
	         : (byte_in == 8'hc8)? 32'hf2c9dd28
	         : (byte_in == 8'hc9)? 32'h476d1b13
	         : (byte_in == 8'hca)? 32'ha1556097
	         : (byte_in == 8'hcb)? 32'h14f1a6ac
	         : (byte_in == 8'hcc)? 32'h7fbc2ad9
	         : (byte_in == 8'hcd)? 32'hca18ece2
	         : (byte_in == 8'hce)? 32'h2c209766
	         : (byte_in == 8'hcf)? 32'h9984515d
	         : (byte_in == 8'hd0)? 32'h4f1b49b4
	         : (byte_in == 8'hd1)? 32'hfabf8f8f
	         : (byte_in == 8'hd2)? 32'h1c87f40b
	         : (byte_in == 8'hd3)? 32'ha9233230
	         : (byte_in == 8'hd4)? 32'hc26ebe45
	         : (byte_in == 8'hd5)? 32'h77ca787e
	         : (byte_in == 8'hd6)? 32'h91f203fa
	         : (byte_in == 8'hd7)? 32'h2456c5c1
	         : (byte_in == 8'hd8)? 32'h5d83f4f2
	         : (byte_in == 8'hd9)? 32'he82732c9
	         : (byte_in == 8'hda)? 32'h0e1f494d
	         : (byte_in == 8'hdb)? 32'hbbbb8f76
	         : (byte_in == 8'hdc)? 32'hd0f60303
	         : (byte_in == 8'hdd)? 32'h6552c538
	         : (byte_in == 8'hde)? 32'h836abebc
	         : (byte_in == 8'hdf)? 32'h36ce7887
	         : (byte_in == 8'he0)? 32'h96fda75d
	         : (byte_in == 8'he1)? 32'h23596166
	         : (byte_in == 8'he2)? 32'hc5611ae2
	         : (byte_in == 8'he3)? 32'h70c5dcd9
	         : (byte_in == 8'he4)? 32'h1b8850ac
	         : (byte_in == 8'he5)? 32'hae2c9697
	         : (byte_in == 8'he6)? 32'h4814ed13
	         : (byte_in == 8'he7)? 32'hfdb02b28
	         : (byte_in == 8'he8)? 32'h84651a1b
	         : (byte_in == 8'he9)? 32'h31c1dc20
	         : (byte_in == 8'hea)? 32'hd7f9a7a4
	         : (byte_in == 8'heb)? 32'h625d619f
	         : (byte_in == 8'hec)? 32'h0910edea
	         : (byte_in == 8'hed)? 32'hbcb42bd1
	         : (byte_in == 8'hee)? 32'h5a8c5055
	         : (byte_in == 8'hef)? 32'hef28966e
	         : (byte_in == 8'hf0)? 32'h39b78e87
	         : (byte_in == 8'hf1)? 32'h8c1348bc
	         : (byte_in == 8'hf2)? 32'h6a2b3338
	         : (byte_in == 8'hf3)? 32'hdf8ff503
	         : (byte_in == 8'hf4)? 32'hb4c27976
	         : (byte_in == 8'hf5)? 32'h0166bf4d
	         : (byte_in == 8'hf6)? 32'he75ec4c9
	         : (byte_in == 8'hf7)? 32'h52fa02f2
	         : (byte_in == 8'hf8)? 32'h2b2f33c1
	         : (byte_in == 8'hf9)? 32'h9e8bf5fa
	         : (byte_in == 8'hfa)? 32'h78b38e7e
	         : (byte_in == 8'hfb)? 32'hcd174845
	         : (byte_in == 8'hfc)? 32'ha65ac430
	         : (byte_in == 8'hfd)? 32'h13fe020b
	         : (byte_in == 8'hfe)? 32'hf5c6798f
	         :                     32'h4062bfb4;

endmodule
//}}}

module TABLE13(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h71575061
	         : (byte_in == 8'h02)? 32'hb1f490bc
	         : (byte_in == 8'h03)? 32'hc0a3c0dd
	         : (byte_in == 8'h04)? 32'he2afa0c0
	         : (byte_in == 8'h05)? 32'h93f8f0a1
	         : (byte_in == 8'h06)? 32'h535b307c
	         : (byte_in == 8'h07)? 32'h220c601d
	         : (byte_in == 8'h08)? 32'h63e92178
	         : (byte_in == 8'h09)? 32'h12be7119
	         : (byte_in == 8'h0a)? 32'hd21db1c4
	         : (byte_in == 8'h0b)? 32'ha34ae1a5
	         : (byte_in == 8'h0c)? 32'h814681b8
	         : (byte_in == 8'h0d)? 32'hf011d1d9
	         : (byte_in == 8'h0e)? 32'h30b21104
	         : (byte_in == 8'h0f)? 32'h41e54165
	         : (byte_in == 8'h10)? 32'h23633a05
	         : (byte_in == 8'h11)? 32'h52346a64
	         : (byte_in == 8'h12)? 32'h9297aab9
	         : (byte_in == 8'h13)? 32'he3c0fad8
	         : (byte_in == 8'h14)? 32'hc1cc9ac5
	         : (byte_in == 8'h15)? 32'hb09bcaa4
	         : (byte_in == 8'h16)? 32'h70380a79
	         : (byte_in == 8'h17)? 32'h016f5a18
	         : (byte_in == 8'h18)? 32'h408a1b7d
	         : (byte_in == 8'h19)? 32'h31dd4b1c
	         : (byte_in == 8'h1a)? 32'hf17e8bc1
	         : (byte_in == 8'h1b)? 32'h8029dba0
	         : (byte_in == 8'h1c)? 32'ha225bbbd
	         : (byte_in == 8'h1d)? 32'hd372ebdc
	         : (byte_in == 8'h1e)? 32'h13d12b01
	         : (byte_in == 8'h1f)? 32'h62867b60
	         : (byte_in == 8'h20)? 32'h727784cb
	         : (byte_in == 8'h21)? 32'h0320d4aa
	         : (byte_in == 8'h22)? 32'hc3831477
	         : (byte_in == 8'h23)? 32'hb2d44416
	         : (byte_in == 8'h24)? 32'h90d8240b
	         : (byte_in == 8'h25)? 32'he18f746a
	         : (byte_in == 8'h26)? 32'h212cb4b7
	         : (byte_in == 8'h27)? 32'h507be4d6
	         : (byte_in == 8'h28)? 32'h119ea5b3
	         : (byte_in == 8'h29)? 32'h60c9f5d2
	         : (byte_in == 8'h2a)? 32'ha06a350f
	         : (byte_in == 8'h2b)? 32'hd13d656e
	         : (byte_in == 8'h2c)? 32'hf3310573
	         : (byte_in == 8'h2d)? 32'h82665512
	         : (byte_in == 8'h2e)? 32'h42c595cf
	         : (byte_in == 8'h2f)? 32'h3392c5ae
	         : (byte_in == 8'h30)? 32'h5114bece
	         : (byte_in == 8'h31)? 32'h2043eeaf
	         : (byte_in == 8'h32)? 32'he0e02e72
	         : (byte_in == 8'h33)? 32'h91b77e13
	         : (byte_in == 8'h34)? 32'hb3bb1e0e
	         : (byte_in == 8'h35)? 32'hc2ec4e6f
	         : (byte_in == 8'h36)? 32'h024f8eb2
	         : (byte_in == 8'h37)? 32'h7318ded3
	         : (byte_in == 8'h38)? 32'h32fd9fb6
	         : (byte_in == 8'h39)? 32'h43aacfd7
	         : (byte_in == 8'h3a)? 32'h83090f0a
	         : (byte_in == 8'h3b)? 32'hf25e5f6b
	         : (byte_in == 8'h3c)? 32'hd0523f76
	         : (byte_in == 8'h3d)? 32'ha1056f17
	         : (byte_in == 8'h3e)? 32'h61a6afca
	         : (byte_in == 8'h3f)? 32'h10f1ffab
	         : (byte_in == 8'h40)? 32'hf362b233
	         : (byte_in == 8'h41)? 32'h8235e252
	         : (byte_in == 8'h42)? 32'h4296228f
	         : (byte_in == 8'h43)? 32'h33c172ee
	         : (byte_in == 8'h44)? 32'h11cd12f3
	         : (byte_in == 8'h45)? 32'h609a4292
	         : (byte_in == 8'h46)? 32'ha039824f
	         : (byte_in == 8'h47)? 32'hd16ed22e
	         : (byte_in == 8'h48)? 32'h908b934b
	         : (byte_in == 8'h49)? 32'he1dcc32a
	         : (byte_in == 8'h4a)? 32'h217f03f7
	         : (byte_in == 8'h4b)? 32'h50285396
	         : (byte_in == 8'h4c)? 32'h7224338b
	         : (byte_in == 8'h4d)? 32'h037363ea
	         : (byte_in == 8'h4e)? 32'hc3d0a337
	         : (byte_in == 8'h4f)? 32'hb287f356
	         : (byte_in == 8'h50)? 32'hd0018836
	         : (byte_in == 8'h51)? 32'ha156d857
	         : (byte_in == 8'h52)? 32'h61f5188a
	         : (byte_in == 8'h53)? 32'h10a248eb
	         : (byte_in == 8'h54)? 32'h32ae28f6
	         : (byte_in == 8'h55)? 32'h43f97897
	         : (byte_in == 8'h56)? 32'h835ab84a
	         : (byte_in == 8'h57)? 32'hf20de82b
	         : (byte_in == 8'h58)? 32'hb3e8a94e
	         : (byte_in == 8'h59)? 32'hc2bff92f
	         : (byte_in == 8'h5a)? 32'h021c39f2
	         : (byte_in == 8'h5b)? 32'h734b6993
	         : (byte_in == 8'h5c)? 32'h5147098e
	         : (byte_in == 8'h5d)? 32'h201059ef
	         : (byte_in == 8'h5e)? 32'he0b39932
	         : (byte_in == 8'h5f)? 32'h91e4c953
	         : (byte_in == 8'h60)? 32'h811536f8
	         : (byte_in == 8'h61)? 32'hf0426699
	         : (byte_in == 8'h62)? 32'h30e1a644
	         : (byte_in == 8'h63)? 32'h41b6f625
	         : (byte_in == 8'h64)? 32'h63ba9638
	         : (byte_in == 8'h65)? 32'h12edc659
	         : (byte_in == 8'h66)? 32'hd24e0684
	         : (byte_in == 8'h67)? 32'ha31956e5
	         : (byte_in == 8'h68)? 32'he2fc1780
	         : (byte_in == 8'h69)? 32'h93ab47e1
	         : (byte_in == 8'h6a)? 32'h5308873c
	         : (byte_in == 8'h6b)? 32'h225fd75d
	         : (byte_in == 8'h6c)? 32'h0053b740
	         : (byte_in == 8'h6d)? 32'h7104e721
	         : (byte_in == 8'h6e)? 32'hb1a727fc
	         : (byte_in == 8'h6f)? 32'hc0f0779d
	         : (byte_in == 8'h70)? 32'ha2760cfd
	         : (byte_in == 8'h71)? 32'hd3215c9c
	         : (byte_in == 8'h72)? 32'h13829c41
	         : (byte_in == 8'h73)? 32'h62d5cc20
	         : (byte_in == 8'h74)? 32'h40d9ac3d
	         : (byte_in == 8'h75)? 32'h318efc5c
	         : (byte_in == 8'h76)? 32'hf12d3c81
	         : (byte_in == 8'h77)? 32'h807a6ce0
	         : (byte_in == 8'h78)? 32'hc19f2d85
	         : (byte_in == 8'h79)? 32'hb0c87de4
	         : (byte_in == 8'h7a)? 32'h706bbd39
	         : (byte_in == 8'h7b)? 32'h013ced58
	         : (byte_in == 8'h7c)? 32'h23308d45
	         : (byte_in == 8'h7d)? 32'h5267dd24
	         : (byte_in == 8'h7e)? 32'h92c41df9
	         : (byte_in == 8'h7f)? 32'he3934d98
	         : (byte_in == 8'h80)? 32'hb772b42b
	         : (byte_in == 8'h81)? 32'hc625e44a
	         : (byte_in == 8'h82)? 32'h06862497
	         : (byte_in == 8'h83)? 32'h77d174f6
	         : (byte_in == 8'h84)? 32'h55dd14eb
	         : (byte_in == 8'h85)? 32'h248a448a
	         : (byte_in == 8'h86)? 32'he4298457
	         : (byte_in == 8'h87)? 32'h957ed436
	         : (byte_in == 8'h88)? 32'hd49b9553
	         : (byte_in == 8'h89)? 32'ha5ccc532
	         : (byte_in == 8'h8a)? 32'h656f05ef
	         : (byte_in == 8'h8b)? 32'h1438558e
	         : (byte_in == 8'h8c)? 32'h36343593
	         : (byte_in == 8'h8d)? 32'h476365f2
	         : (byte_in == 8'h8e)? 32'h87c0a52f
	         : (byte_in == 8'h8f)? 32'hf697f54e
	         : (byte_in == 8'h90)? 32'h94118e2e
	         : (byte_in == 8'h91)? 32'he546de4f
	         : (byte_in == 8'h92)? 32'h25e51e92
	         : (byte_in == 8'h93)? 32'h54b24ef3
	         : (byte_in == 8'h94)? 32'h76be2eee
	         : (byte_in == 8'h95)? 32'h07e97e8f
	         : (byte_in == 8'h96)? 32'hc74abe52
	         : (byte_in == 8'h97)? 32'hb61dee33
	         : (byte_in == 8'h98)? 32'hf7f8af56
	         : (byte_in == 8'h99)? 32'h86afff37
	         : (byte_in == 8'h9a)? 32'h460c3fea
	         : (byte_in == 8'h9b)? 32'h375b6f8b
	         : (byte_in == 8'h9c)? 32'h15570f96
	         : (byte_in == 8'h9d)? 32'h64005ff7
	         : (byte_in == 8'h9e)? 32'ha4a39f2a
	         : (byte_in == 8'h9f)? 32'hd5f4cf4b
	         : (byte_in == 8'ha0)? 32'hc50530e0
	         : (byte_in == 8'ha1)? 32'hb4526081
	         : (byte_in == 8'ha2)? 32'h74f1a05c
	         : (byte_in == 8'ha3)? 32'h05a6f03d
	         : (byte_in == 8'ha4)? 32'h27aa9020
	         : (byte_in == 8'ha5)? 32'h56fdc041
	         : (byte_in == 8'ha6)? 32'h965e009c
	         : (byte_in == 8'ha7)? 32'he70950fd
	         : (byte_in == 8'ha8)? 32'ha6ec1198
	         : (byte_in == 8'ha9)? 32'hd7bb41f9
	         : (byte_in == 8'haa)? 32'h17188124
	         : (byte_in == 8'hab)? 32'h664fd145
	         : (byte_in == 8'hac)? 32'h4443b158
	         : (byte_in == 8'had)? 32'h3514e139
	         : (byte_in == 8'hae)? 32'hf5b721e4
	         : (byte_in == 8'haf)? 32'h84e07185
	         : (byte_in == 8'hb0)? 32'he6660ae5
	         : (byte_in == 8'hb1)? 32'h97315a84
	         : (byte_in == 8'hb2)? 32'h57929a59
	         : (byte_in == 8'hb3)? 32'h26c5ca38
	         : (byte_in == 8'hb4)? 32'h04c9aa25
	         : (byte_in == 8'hb5)? 32'h759efa44
	         : (byte_in == 8'hb6)? 32'hb53d3a99
	         : (byte_in == 8'hb7)? 32'hc46a6af8
	         : (byte_in == 8'hb8)? 32'h858f2b9d
	         : (byte_in == 8'hb9)? 32'hf4d87bfc
	         : (byte_in == 8'hba)? 32'h347bbb21
	         : (byte_in == 8'hbb)? 32'h452ceb40
	         : (byte_in == 8'hbc)? 32'h67208b5d
	         : (byte_in == 8'hbd)? 32'h1677db3c
	         : (byte_in == 8'hbe)? 32'hd6d41be1
	         : (byte_in == 8'hbf)? 32'ha7834b80
	         : (byte_in == 8'hc0)? 32'h44100618
	         : (byte_in == 8'hc1)? 32'h35475679
	         : (byte_in == 8'hc2)? 32'hf5e496a4
	         : (byte_in == 8'hc3)? 32'h84b3c6c5
	         : (byte_in == 8'hc4)? 32'ha6bfa6d8
	         : (byte_in == 8'hc5)? 32'hd7e8f6b9
	         : (byte_in == 8'hc6)? 32'h174b3664
	         : (byte_in == 8'hc7)? 32'h661c6605
	         : (byte_in == 8'hc8)? 32'h27f92760
	         : (byte_in == 8'hc9)? 32'h56ae7701
	         : (byte_in == 8'hca)? 32'h960db7dc
	         : (byte_in == 8'hcb)? 32'he75ae7bd
	         : (byte_in == 8'hcc)? 32'hc55687a0
	         : (byte_in == 8'hcd)? 32'hb401d7c1
	         : (byte_in == 8'hce)? 32'h74a2171c
	         : (byte_in == 8'hcf)? 32'h05f5477d
	         : (byte_in == 8'hd0)? 32'h67733c1d
	         : (byte_in == 8'hd1)? 32'h16246c7c
	         : (byte_in == 8'hd2)? 32'hd687aca1
	         : (byte_in == 8'hd3)? 32'ha7d0fcc0
	         : (byte_in == 8'hd4)? 32'h85dc9cdd
	         : (byte_in == 8'hd5)? 32'hf48bccbc
	         : (byte_in == 8'hd6)? 32'h34280c61
	         : (byte_in == 8'hd7)? 32'h457f5c00
	         : (byte_in == 8'hd8)? 32'h049a1d65
	         : (byte_in == 8'hd9)? 32'h75cd4d04
	         : (byte_in == 8'hda)? 32'hb56e8dd9
	         : (byte_in == 8'hdb)? 32'hc439ddb8
	         : (byte_in == 8'hdc)? 32'he635bda5
	         : (byte_in == 8'hdd)? 32'h9762edc4
	         : (byte_in == 8'hde)? 32'h57c12d19
	         : (byte_in == 8'hdf)? 32'h26967d78
	         : (byte_in == 8'he0)? 32'h366782d3
	         : (byte_in == 8'he1)? 32'h4730d2b2
	         : (byte_in == 8'he2)? 32'h8793126f
	         : (byte_in == 8'he3)? 32'hf6c4420e
	         : (byte_in == 8'he4)? 32'hd4c82213
	         : (byte_in == 8'he5)? 32'ha59f7272
	         : (byte_in == 8'he6)? 32'h653cb2af
	         : (byte_in == 8'he7)? 32'h146be2ce
	         : (byte_in == 8'he8)? 32'h558ea3ab
	         : (byte_in == 8'he9)? 32'h24d9f3ca
	         : (byte_in == 8'hea)? 32'he47a3317
	         : (byte_in == 8'heb)? 32'h952d6376
	         : (byte_in == 8'hec)? 32'hb721036b
	         : (byte_in == 8'hed)? 32'hc676530a
	         : (byte_in == 8'hee)? 32'h06d593d7
	         : (byte_in == 8'hef)? 32'h7782c3b6
	         : (byte_in == 8'hf0)? 32'h1504b8d6
	         : (byte_in == 8'hf1)? 32'h6453e8b7
	         : (byte_in == 8'hf2)? 32'ha4f0286a
	         : (byte_in == 8'hf3)? 32'hd5a7780b
	         : (byte_in == 8'hf4)? 32'hf7ab1816
	         : (byte_in == 8'hf5)? 32'h86fc4877
	         : (byte_in == 8'hf6)? 32'h465f88aa
	         : (byte_in == 8'hf7)? 32'h3708d8cb
	         : (byte_in == 8'hf8)? 32'h76ed99ae
	         : (byte_in == 8'hf9)? 32'h07bac9cf
	         : (byte_in == 8'hfa)? 32'hc7190912
	         : (byte_in == 8'hfb)? 32'hb64e5973
	         : (byte_in == 8'hfc)? 32'h9442396e
	         : (byte_in == 8'hfd)? 32'he515690f
	         : (byte_in == 8'hfe)? 32'h25b6a9d2
	         :                     32'h54e1f9b3;

endmodule
//}}}

module TABLE14(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'he6c46464
	         : (byte_in == 8'h02)? 32'h6ee56854
	         : (byte_in == 8'h03)? 32'h88210c30
	         : (byte_in == 8'h04)? 32'h9e147576
	         : (byte_in == 8'h05)? 32'h78d01112
	         : (byte_in == 8'h06)? 32'hf0f11d22
	         : (byte_in == 8'h07)? 32'h16357946
	         : (byte_in == 8'h08)? 32'h3bf3ab2c
	         : (byte_in == 8'h09)? 32'hdd37cf48
	         : (byte_in == 8'h0a)? 32'h5516c378
	         : (byte_in == 8'h0b)? 32'hb3d2a71c
	         : (byte_in == 8'h0c)? 32'ha5e7de5a
	         : (byte_in == 8'h0d)? 32'h4323ba3e
	         : (byte_in == 8'h0e)? 32'hcb02b60e
	         : (byte_in == 8'h0f)? 32'h2dc6d26a
	         : (byte_in == 8'h10)? 32'h898d2cd6
	         : (byte_in == 8'h11)? 32'h6f4948b2
	         : (byte_in == 8'h12)? 32'he7684482
	         : (byte_in == 8'h13)? 32'h01ac20e6
	         : (byte_in == 8'h14)? 32'h179959a0
	         : (byte_in == 8'h15)? 32'hf15d3dc4
	         : (byte_in == 8'h16)? 32'h797c31f4
	         : (byte_in == 8'h17)? 32'h9fb85590
	         : (byte_in == 8'h18)? 32'hb27e87fa
	         : (byte_in == 8'h19)? 32'h54bae39e
	         : (byte_in == 8'h1a)? 32'hdc9befae
	         : (byte_in == 8'h1b)? 32'h3a5f8bca
	         : (byte_in == 8'h1c)? 32'h2c6af28c
	         : (byte_in == 8'h1d)? 32'hcaae96e8
	         : (byte_in == 8'h1e)? 32'h428f9ad8
	         : (byte_in == 8'h1f)? 32'ha44bfebc
	         : (byte_in == 8'h20)? 32'h247febe6
	         : (byte_in == 8'h21)? 32'hc2bb8f82
	         : (byte_in == 8'h22)? 32'h4a9a83b2
	         : (byte_in == 8'h23)? 32'hac5ee7d6
	         : (byte_in == 8'h24)? 32'hba6b9e90
	         : (byte_in == 8'h25)? 32'h5caffaf4
	         : (byte_in == 8'h26)? 32'hd48ef6c4
	         : (byte_in == 8'h27)? 32'h324a92a0
	         : (byte_in == 8'h28)? 32'h1f8c40ca
	         : (byte_in == 8'h29)? 32'hf94824ae
	         : (byte_in == 8'h2a)? 32'h7169289e
	         : (byte_in == 8'h2b)? 32'h97ad4cfa
	         : (byte_in == 8'h2c)? 32'h819835bc
	         : (byte_in == 8'h2d)? 32'h675c51d8
	         : (byte_in == 8'h2e)? 32'hef7d5de8
	         : (byte_in == 8'h2f)? 32'h09b9398c
	         : (byte_in == 8'h30)? 32'hadf2c730
	         : (byte_in == 8'h31)? 32'h4b36a354
	         : (byte_in == 8'h32)? 32'hc317af64
	         : (byte_in == 8'h33)? 32'h25d3cb00
	         : (byte_in == 8'h34)? 32'h33e6b246
	         : (byte_in == 8'h35)? 32'hd522d622
	         : (byte_in == 8'h36)? 32'h5d03da12
	         : (byte_in == 8'h37)? 32'hbbc7be76
	         : (byte_in == 8'h38)? 32'h96016c1c
	         : (byte_in == 8'h39)? 32'h70c50878
	         : (byte_in == 8'h3a)? 32'hf8e40448
	         : (byte_in == 8'h3b)? 32'h1e20602c
	         : (byte_in == 8'h3c)? 32'h0815196a
	         : (byte_in == 8'h3d)? 32'heed17d0e
	         : (byte_in == 8'h3e)? 32'h66f0713e
	         : (byte_in == 8'h3f)? 32'h8034155a
	         : (byte_in == 8'h40)? 32'ha6bf9f96
	         : (byte_in == 8'h41)? 32'h407bfbf2
	         : (byte_in == 8'h42)? 32'hc85af7c2
	         : (byte_in == 8'h43)? 32'h2e9e93a6
	         : (byte_in == 8'h44)? 32'h38abeae0
	         : (byte_in == 8'h45)? 32'hde6f8e84
	         : (byte_in == 8'h46)? 32'h564e82b4
	         : (byte_in == 8'h47)? 32'hb08ae6d0
	         : (byte_in == 8'h48)? 32'h9d4c34ba
	         : (byte_in == 8'h49)? 32'h7b8850de
	         : (byte_in == 8'h4a)? 32'hf3a95cee
	         : (byte_in == 8'h4b)? 32'h156d388a
	         : (byte_in == 8'h4c)? 32'h035841cc
	         : (byte_in == 8'h4d)? 32'he59c25a8
	         : (byte_in == 8'h4e)? 32'h6dbd2998
	         : (byte_in == 8'h4f)? 32'h8b794dfc
	         : (byte_in == 8'h50)? 32'h2f32b340
	         : (byte_in == 8'h51)? 32'hc9f6d724
	         : (byte_in == 8'h52)? 32'h41d7db14
	         : (byte_in == 8'h53)? 32'ha713bf70
	         : (byte_in == 8'h54)? 32'hb126c636
	         : (byte_in == 8'h55)? 32'h57e2a252
	         : (byte_in == 8'h56)? 32'hdfc3ae62
	         : (byte_in == 8'h57)? 32'h3907ca06
	         : (byte_in == 8'h58)? 32'h14c1186c
	         : (byte_in == 8'h59)? 32'hf2057c08
	         : (byte_in == 8'h5a)? 32'h7a247038
	         : (byte_in == 8'h5b)? 32'h9ce0145c
	         : (byte_in == 8'h5c)? 32'h8ad56d1a
	         : (byte_in == 8'h5d)? 32'h6c11097e
	         : (byte_in == 8'h5e)? 32'he430054e
	         : (byte_in == 8'h5f)? 32'h02f4612a
	         : (byte_in == 8'h60)? 32'h82c07470
	         : (byte_in == 8'h61)? 32'h64041014
	         : (byte_in == 8'h62)? 32'hec251c24
	         : (byte_in == 8'h63)? 32'h0ae17840
	         : (byte_in == 8'h64)? 32'h1cd40106
	         : (byte_in == 8'h65)? 32'hfa106562
	         : (byte_in == 8'h66)? 32'h72316952
	         : (byte_in == 8'h67)? 32'h94f50d36
	         : (byte_in == 8'h68)? 32'hb933df5c
	         : (byte_in == 8'h69)? 32'h5ff7bb38
	         : (byte_in == 8'h6a)? 32'hd7d6b708
	         : (byte_in == 8'h6b)? 32'h3112d36c
	         : (byte_in == 8'h6c)? 32'h2727aa2a
	         : (byte_in == 8'h6d)? 32'hc1e3ce4e
	         : (byte_in == 8'h6e)? 32'h49c2c27e
	         : (byte_in == 8'h6f)? 32'haf06a61a
	         : (byte_in == 8'h70)? 32'h0b4d58a6
	         : (byte_in == 8'h71)? 32'hed893cc2
	         : (byte_in == 8'h72)? 32'h65a830f2
	         : (byte_in == 8'h73)? 32'h836c5496
	         : (byte_in == 8'h74)? 32'h95592dd0
	         : (byte_in == 8'h75)? 32'h739d49b4
	         : (byte_in == 8'h76)? 32'hfbbc4584
	         : (byte_in == 8'h77)? 32'h1d7821e0
	         : (byte_in == 8'h78)? 32'h30bef38a
	         : (byte_in == 8'h79)? 32'hd67a97ee
	         : (byte_in == 8'h7a)? 32'h5e5b9bde
	         : (byte_in == 8'h7b)? 32'hb89fffba
	         : (byte_in == 8'h7c)? 32'haeaa86fc
	         : (byte_in == 8'h7d)? 32'h486ee298
	         : (byte_in == 8'h7e)? 32'hc04feea8
	         : (byte_in == 8'h7f)? 32'h268b8acc
	         : (byte_in == 8'h80)? 32'h1b666a73
	         : (byte_in == 8'h81)? 32'hfda20e17
	         : (byte_in == 8'h82)? 32'h75830227
	         : (byte_in == 8'h83)? 32'h93476643
	         : (byte_in == 8'h84)? 32'h85721f05
	         : (byte_in == 8'h85)? 32'h63b67b61
	         : (byte_in == 8'h86)? 32'heb977751
	         : (byte_in == 8'h87)? 32'h0d531335
	         : (byte_in == 8'h88)? 32'h2095c15f
	         : (byte_in == 8'h89)? 32'hc651a53b
	         : (byte_in == 8'h8a)? 32'h4e70a90b
	         : (byte_in == 8'h8b)? 32'ha8b4cd6f
	         : (byte_in == 8'h8c)? 32'hbe81b429
	         : (byte_in == 8'h8d)? 32'h5845d04d
	         : (byte_in == 8'h8e)? 32'hd064dc7d
	         : (byte_in == 8'h8f)? 32'h36a0b819
	         : (byte_in == 8'h90)? 32'h92eb46a5
	         : (byte_in == 8'h91)? 32'h742f22c1
	         : (byte_in == 8'h92)? 32'hfc0e2ef1
	         : (byte_in == 8'h93)? 32'h1aca4a95
	         : (byte_in == 8'h94)? 32'h0cff33d3
	         : (byte_in == 8'h95)? 32'hea3b57b7
	         : (byte_in == 8'h96)? 32'h621a5b87
	         : (byte_in == 8'h97)? 32'h84de3fe3
	         : (byte_in == 8'h98)? 32'ha918ed89
	         : (byte_in == 8'h99)? 32'h4fdc89ed
	         : (byte_in == 8'h9a)? 32'hc7fd85dd
	         : (byte_in == 8'h9b)? 32'h2139e1b9
	         : (byte_in == 8'h9c)? 32'h370c98ff
	         : (byte_in == 8'h9d)? 32'hd1c8fc9b
	         : (byte_in == 8'h9e)? 32'h59e9f0ab
	         : (byte_in == 8'h9f)? 32'hbf2d94cf
	         : (byte_in == 8'ha0)? 32'h3f198195
	         : (byte_in == 8'ha1)? 32'hd9dde5f1
	         : (byte_in == 8'ha2)? 32'h51fce9c1
	         : (byte_in == 8'ha3)? 32'hb7388da5
	         : (byte_in == 8'ha4)? 32'ha10df4e3
	         : (byte_in == 8'ha5)? 32'h47c99087
	         : (byte_in == 8'ha6)? 32'hcfe89cb7
	         : (byte_in == 8'ha7)? 32'h292cf8d3
	         : (byte_in == 8'ha8)? 32'h04ea2ab9
	         : (byte_in == 8'ha9)? 32'he22e4edd
	         : (byte_in == 8'haa)? 32'h6a0f42ed
	         : (byte_in == 8'hab)? 32'h8ccb2689
	         : (byte_in == 8'hac)? 32'h9afe5fcf
	         : (byte_in == 8'had)? 32'h7c3a3bab
	         : (byte_in == 8'hae)? 32'hf41b379b
	         : (byte_in == 8'haf)? 32'h12df53ff
	         : (byte_in == 8'hb0)? 32'hb694ad43
	         : (byte_in == 8'hb1)? 32'h5050c927
	         : (byte_in == 8'hb2)? 32'hd871c517
	         : (byte_in == 8'hb3)? 32'h3eb5a173
	         : (byte_in == 8'hb4)? 32'h2880d835
	         : (byte_in == 8'hb5)? 32'hce44bc51
	         : (byte_in == 8'hb6)? 32'h4665b061
	         : (byte_in == 8'hb7)? 32'ha0a1d405
	         : (byte_in == 8'hb8)? 32'h8d67066f
	         : (byte_in == 8'hb9)? 32'h6ba3620b
	         : (byte_in == 8'hba)? 32'he3826e3b
	         : (byte_in == 8'hbb)? 32'h05460a5f
	         : (byte_in == 8'hbc)? 32'h13737319
	         : (byte_in == 8'hbd)? 32'hf5b7177d
	         : (byte_in == 8'hbe)? 32'h7d961b4d
	         : (byte_in == 8'hbf)? 32'h9b527f29
	         : (byte_in == 8'hc0)? 32'hbdd9f5e5
	         : (byte_in == 8'hc1)? 32'h5b1d9181
	         : (byte_in == 8'hc2)? 32'hd33c9db1
	         : (byte_in == 8'hc3)? 32'h35f8f9d5
	         : (byte_in == 8'hc4)? 32'h23cd8093
	         : (byte_in == 8'hc5)? 32'hc509e4f7
	         : (byte_in == 8'hc6)? 32'h4d28e8c7
	         : (byte_in == 8'hc7)? 32'habec8ca3
	         : (byte_in == 8'hc8)? 32'h862a5ec9
	         : (byte_in == 8'hc9)? 32'h60ee3aad
	         : (byte_in == 8'hca)? 32'he8cf369d
	         : (byte_in == 8'hcb)? 32'h0e0b52f9
	         : (byte_in == 8'hcc)? 32'h183e2bbf
	         : (byte_in == 8'hcd)? 32'hfefa4fdb
	         : (byte_in == 8'hce)? 32'h76db43eb
	         : (byte_in == 8'hcf)? 32'h901f278f
	         : (byte_in == 8'hd0)? 32'h3454d933
	         : (byte_in == 8'hd1)? 32'hd290bd57
	         : (byte_in == 8'hd2)? 32'h5ab1b167
	         : (byte_in == 8'hd3)? 32'hbc75d503
	         : (byte_in == 8'hd4)? 32'haa40ac45
	         : (byte_in == 8'hd5)? 32'h4c84c821
	         : (byte_in == 8'hd6)? 32'hc4a5c411
	         : (byte_in == 8'hd7)? 32'h2261a075
	         : (byte_in == 8'hd8)? 32'h0fa7721f
	         : (byte_in == 8'hd9)? 32'he963167b
	         : (byte_in == 8'hda)? 32'h61421a4b
	         : (byte_in == 8'hdb)? 32'h87867e2f
	         : (byte_in == 8'hdc)? 32'h91b30769
	         : (byte_in == 8'hdd)? 32'h7777630d
	         : (byte_in == 8'hde)? 32'hff566f3d
	         : (byte_in == 8'hdf)? 32'h19920b59
	         : (byte_in == 8'he0)? 32'h99a61e03
	         : (byte_in == 8'he1)? 32'h7f627a67
	         : (byte_in == 8'he2)? 32'hf7437657
	         : (byte_in == 8'he3)? 32'h11871233
	         : (byte_in == 8'he4)? 32'h07b26b75
	         : (byte_in == 8'he5)? 32'he1760f11
	         : (byte_in == 8'he6)? 32'h69570321
	         : (byte_in == 8'he7)? 32'h8f936745
	         : (byte_in == 8'he8)? 32'ha255b52f
	         : (byte_in == 8'he9)? 32'h4491d14b
	         : (byte_in == 8'hea)? 32'hccb0dd7b
	         : (byte_in == 8'heb)? 32'h2a74b91f
	         : (byte_in == 8'hec)? 32'h3c41c059
	         : (byte_in == 8'hed)? 32'hda85a43d
	         : (byte_in == 8'hee)? 32'h52a4a80d
	         : (byte_in == 8'hef)? 32'hb460cc69
	         : (byte_in == 8'hf0)? 32'h102b32d5
	         : (byte_in == 8'hf1)? 32'hf6ef56b1
	         : (byte_in == 8'hf2)? 32'h7ece5a81
	         : (byte_in == 8'hf3)? 32'h980a3ee5
	         : (byte_in == 8'hf4)? 32'h8e3f47a3
	         : (byte_in == 8'hf5)? 32'h68fb23c7
	         : (byte_in == 8'hf6)? 32'he0da2ff7
	         : (byte_in == 8'hf7)? 32'h061e4b93
	         : (byte_in == 8'hf8)? 32'h2bd899f9
	         : (byte_in == 8'hf9)? 32'hcd1cfd9d
	         : (byte_in == 8'hfa)? 32'h453df1ad
	         : (byte_in == 8'hfb)? 32'ha3f995c9
	         : (byte_in == 8'hfc)? 32'hb5ccec8f
	         : (byte_in == 8'hfd)? 32'h530888eb
	         : (byte_in == 8'hfe)? 32'hdb2984db
	         :                     32'h3dede0bf;

endmodule
//}}}

module TABLE15(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h1ee68292
	         : (byte_in == 8'h02)? 32'hd0f4af61
	         : (byte_in == 8'h03)? 32'hce122df3
	         : (byte_in == 8'h04)? 32'h3dc90524
	         : (byte_in == 8'h05)? 32'h232f87b6
	         : (byte_in == 8'h06)? 32'hed3daa45
	         : (byte_in == 8'h07)? 32'hf3db28d7
	         : (byte_in == 8'h08)? 32'ha1ec5ec1
	         : (byte_in == 8'h09)? 32'hbf0adc53
	         : (byte_in == 8'h0a)? 32'h7118f1a0
	         : (byte_in == 8'h0b)? 32'h6ffe7332
	         : (byte_in == 8'h0c)? 32'h9c255be5
	         : (byte_in == 8'h0d)? 32'h82c3d977
	         : (byte_in == 8'h0e)? 32'h4cd1f484
	         : (byte_in == 8'h0f)? 32'h52377616
	         : (byte_in == 8'h10)? 32'hce36cc72
	         : (byte_in == 8'h11)? 32'hd0d04ee0
	         : (byte_in == 8'h12)? 32'h1ec26313
	         : (byte_in == 8'h13)? 32'h0024e181
	         : (byte_in == 8'h14)? 32'hf3ffc956
	         : (byte_in == 8'h15)? 32'hed194bc4
	         : (byte_in == 8'h16)? 32'h230b6637
	         : (byte_in == 8'h17)? 32'h3dede4a5
	         : (byte_in == 8'h18)? 32'h6fda92b3
	         : (byte_in == 8'h19)? 32'h713c1021
	         : (byte_in == 8'h1a)? 32'hbf2e3dd2
	         : (byte_in == 8'h1b)? 32'ha1c8bf40
	         : (byte_in == 8'h1c)? 32'h52139797
	         : (byte_in == 8'h1d)? 32'h4cf51505
	         : (byte_in == 8'h1e)? 32'h82e738f6
	         : (byte_in == 8'h1f)? 32'h9c01ba64
	         : (byte_in == 8'h20)? 32'h1041003e
	         : (byte_in == 8'h21)? 32'h0ea782ac
	         : (byte_in == 8'h22)? 32'hc0b5af5f
	         : (byte_in == 8'h23)? 32'hde532dcd
	         : (byte_in == 8'h24)? 32'h2d88051a
	         : (byte_in == 8'h25)? 32'h336e8788
	         : (byte_in == 8'h26)? 32'hfd7caa7b
	         : (byte_in == 8'h27)? 32'he39a28e9
	         : (byte_in == 8'h28)? 32'hb1ad5eff
	         : (byte_in == 8'h29)? 32'haf4bdc6d
	         : (byte_in == 8'h2a)? 32'h6159f19e
	         : (byte_in == 8'h2b)? 32'h7fbf730c
	         : (byte_in == 8'h2c)? 32'h8c645bdb
	         : (byte_in == 8'h2d)? 32'h9282d949
	         : (byte_in == 8'h2e)? 32'h5c90f4ba
	         : (byte_in == 8'h2f)? 32'h42767628
	         : (byte_in == 8'h30)? 32'hde77cc4c
	         : (byte_in == 8'h31)? 32'hc0914ede
	         : (byte_in == 8'h32)? 32'h0e83632d
	         : (byte_in == 8'h33)? 32'h1065e1bf
	         : (byte_in == 8'h34)? 32'he3bec968
	         : (byte_in == 8'h35)? 32'hfd584bfa
	         : (byte_in == 8'h36)? 32'h334a6609
	         : (byte_in == 8'h37)? 32'h2dace49b
	         : (byte_in == 8'h38)? 32'h7f9b928d
	         : (byte_in == 8'h39)? 32'h617d101f
	         : (byte_in == 8'h3a)? 32'haf6f3dec
	         : (byte_in == 8'h3b)? 32'hb189bf7e
	         : (byte_in == 8'h3c)? 32'h425297a9
	         : (byte_in == 8'h3d)? 32'h5cb4153b
	         : (byte_in == 8'h3e)? 32'h92a638c8
	         : (byte_in == 8'h3f)? 32'h8c40ba5a
	         : (byte_in == 8'h40)? 32'h29cc5edf
	         : (byte_in == 8'h41)? 32'h372adc4d
	         : (byte_in == 8'h42)? 32'hf938f1be
	         : (byte_in == 8'h43)? 32'he7de732c
	         : (byte_in == 8'h44)? 32'h14055bfb
	         : (byte_in == 8'h45)? 32'h0ae3d969
	         : (byte_in == 8'h46)? 32'hc4f1f49a
	         : (byte_in == 8'h47)? 32'hda177608
	         : (byte_in == 8'h48)? 32'h8820001e
	         : (byte_in == 8'h49)? 32'h96c6828c
	         : (byte_in == 8'h4a)? 32'h58d4af7f
	         : (byte_in == 8'h4b)? 32'h46322ded
	         : (byte_in == 8'h4c)? 32'hb5e9053a
	         : (byte_in == 8'h4d)? 32'hab0f87a8
	         : (byte_in == 8'h4e)? 32'h651daa5b
	         : (byte_in == 8'h4f)? 32'h7bfb28c9
	         : (byte_in == 8'h50)? 32'he7fa92ad
	         : (byte_in == 8'h51)? 32'hf91c103f
	         : (byte_in == 8'h52)? 32'h370e3dcc
	         : (byte_in == 8'h53)? 32'h29e8bf5e
	         : (byte_in == 8'h54)? 32'hda339789
	         : (byte_in == 8'h55)? 32'hc4d5151b
	         : (byte_in == 8'h56)? 32'h0ac738e8
	         : (byte_in == 8'h57)? 32'h1421ba7a
	         : (byte_in == 8'h58)? 32'h4616cc6c
	         : (byte_in == 8'h59)? 32'h58f04efe
	         : (byte_in == 8'h5a)? 32'h96e2630d
	         : (byte_in == 8'h5b)? 32'h8804e19f
	         : (byte_in == 8'h5c)? 32'h7bdfc948
	         : (byte_in == 8'h5d)? 32'h65394bda
	         : (byte_in == 8'h5e)? 32'hab2b6629
	         : (byte_in == 8'h5f)? 32'hb5cde4bb
	         : (byte_in == 8'h60)? 32'h398d5ee1
	         : (byte_in == 8'h61)? 32'h276bdc73
	         : (byte_in == 8'h62)? 32'he979f180
	         : (byte_in == 8'h63)? 32'hf79f7312
	         : (byte_in == 8'h64)? 32'h04445bc5
	         : (byte_in == 8'h65)? 32'h1aa2d957
	         : (byte_in == 8'h66)? 32'hd4b0f4a4
	         : (byte_in == 8'h67)? 32'hca567636
	         : (byte_in == 8'h68)? 32'h98610020
	         : (byte_in == 8'h69)? 32'h868782b2
	         : (byte_in == 8'h6a)? 32'h4895af41
	         : (byte_in == 8'h6b)? 32'h56732dd3
	         : (byte_in == 8'h6c)? 32'ha5a80504
	         : (byte_in == 8'h6d)? 32'hbb4e8796
	         : (byte_in == 8'h6e)? 32'h755caa65
	         : (byte_in == 8'h6f)? 32'h6bba28f7
	         : (byte_in == 8'h70)? 32'hf7bb9293
	         : (byte_in == 8'h71)? 32'he95d1001
	         : (byte_in == 8'h72)? 32'h274f3df2
	         : (byte_in == 8'h73)? 32'h39a9bf60
	         : (byte_in == 8'h74)? 32'hca7297b7
	         : (byte_in == 8'h75)? 32'hd4941525
	         : (byte_in == 8'h76)? 32'h1a8638d6
	         : (byte_in == 8'h77)? 32'h0460ba44
	         : (byte_in == 8'h78)? 32'h5657cc52
	         : (byte_in == 8'h79)? 32'h48b14ec0
	         : (byte_in == 8'h7a)? 32'h86a36333
	         : (byte_in == 8'h7b)? 32'h9845e1a1
	         : (byte_in == 8'h7c)? 32'h6b9ec976
	         : (byte_in == 8'h7d)? 32'h75784be4
	         : (byte_in == 8'h7e)? 32'hbb6a6617
	         : (byte_in == 8'h7f)? 32'ha58ce485
	         : (byte_in == 8'h80)? 32'h731ebdc2
	         : (byte_in == 8'h81)? 32'h6df83f50
	         : (byte_in == 8'h82)? 32'ha3ea12a3
	         : (byte_in == 8'h83)? 32'hbd0c9031
	         : (byte_in == 8'h84)? 32'h4ed7b8e6
	         : (byte_in == 8'h85)? 32'h50313a74
	         : (byte_in == 8'h86)? 32'h9e231787
	         : (byte_in == 8'h87)? 32'h80c59515
	         : (byte_in == 8'h88)? 32'hd2f2e303
	         : (byte_in == 8'h89)? 32'hcc146191
	         : (byte_in == 8'h8a)? 32'h02064c62
	         : (byte_in == 8'h8b)? 32'h1ce0cef0
	         : (byte_in == 8'h8c)? 32'hef3be627
	         : (byte_in == 8'h8d)? 32'hf1dd64b5
	         : (byte_in == 8'h8e)? 32'h3fcf4946
	         : (byte_in == 8'h8f)? 32'h2129cbd4
	         : (byte_in == 8'h90)? 32'hbd2871b0
	         : (byte_in == 8'h91)? 32'ha3cef322
	         : (byte_in == 8'h92)? 32'h6ddcded1
	         : (byte_in == 8'h93)? 32'h733a5c43
	         : (byte_in == 8'h94)? 32'h80e17494
	         : (byte_in == 8'h95)? 32'h9e07f606
	         : (byte_in == 8'h96)? 32'h5015dbf5
	         : (byte_in == 8'h97)? 32'h4ef35967
	         : (byte_in == 8'h98)? 32'h1cc42f71
	         : (byte_in == 8'h99)? 32'h0222ade3
	         : (byte_in == 8'h9a)? 32'hcc308010
	         : (byte_in == 8'h9b)? 32'hd2d60282
	         : (byte_in == 8'h9c)? 32'h210d2a55
	         : (byte_in == 8'h9d)? 32'h3feba8c7
	         : (byte_in == 8'h9e)? 32'hf1f98534
	         : (byte_in == 8'h9f)? 32'hef1f07a6
	         : (byte_in == 8'ha0)? 32'h635fbdfc
	         : (byte_in == 8'ha1)? 32'h7db93f6e
	         : (byte_in == 8'ha2)? 32'hb3ab129d
	         : (byte_in == 8'ha3)? 32'had4d900f
	         : (byte_in == 8'ha4)? 32'h5e96b8d8
	         : (byte_in == 8'ha5)? 32'h40703a4a
	         : (byte_in == 8'ha6)? 32'h8e6217b9
	         : (byte_in == 8'ha7)? 32'h9084952b
	         : (byte_in == 8'ha8)? 32'hc2b3e33d
	         : (byte_in == 8'ha9)? 32'hdc5561af
	         : (byte_in == 8'haa)? 32'h12474c5c
	         : (byte_in == 8'hab)? 32'h0ca1cece
	         : (byte_in == 8'hac)? 32'hff7ae619
	         : (byte_in == 8'had)? 32'he19c648b
	         : (byte_in == 8'hae)? 32'h2f8e4978
	         : (byte_in == 8'haf)? 32'h3168cbea
	         : (byte_in == 8'hb0)? 32'had69718e
	         : (byte_in == 8'hb1)? 32'hb38ff31c
	         : (byte_in == 8'hb2)? 32'h7d9ddeef
	         : (byte_in == 8'hb3)? 32'h637b5c7d
	         : (byte_in == 8'hb4)? 32'h90a074aa
	         : (byte_in == 8'hb5)? 32'h8e46f638
	         : (byte_in == 8'hb6)? 32'h4054dbcb
	         : (byte_in == 8'hb7)? 32'h5eb25959
	         : (byte_in == 8'hb8)? 32'h0c852f4f
	         : (byte_in == 8'hb9)? 32'h1263addd
	         : (byte_in == 8'hba)? 32'hdc71802e
	         : (byte_in == 8'hbb)? 32'hc29702bc
	         : (byte_in == 8'hbc)? 32'h314c2a6b
	         : (byte_in == 8'hbd)? 32'h2faaa8f9
	         : (byte_in == 8'hbe)? 32'he1b8850a
	         : (byte_in == 8'hbf)? 32'hff5e0798
	         : (byte_in == 8'hc0)? 32'h5ad2e31d
	         : (byte_in == 8'hc1)? 32'h4434618f
	         : (byte_in == 8'hc2)? 32'h8a264c7c
	         : (byte_in == 8'hc3)? 32'h94c0ceee
	         : (byte_in == 8'hc4)? 32'h671be639
	         : (byte_in == 8'hc5)? 32'h79fd64ab
	         : (byte_in == 8'hc6)? 32'hb7ef4958
	         : (byte_in == 8'hc7)? 32'ha909cbca
	         : (byte_in == 8'hc8)? 32'hfb3ebddc
	         : (byte_in == 8'hc9)? 32'he5d83f4e
	         : (byte_in == 8'hca)? 32'h2bca12bd
	         : (byte_in == 8'hcb)? 32'h352c902f
	         : (byte_in == 8'hcc)? 32'hc6f7b8f8
	         : (byte_in == 8'hcd)? 32'hd8113a6a
	         : (byte_in == 8'hce)? 32'h16031799
	         : (byte_in == 8'hcf)? 32'h08e5950b
	         : (byte_in == 8'hd0)? 32'h94e42f6f
	         : (byte_in == 8'hd1)? 32'h8a02adfd
	         : (byte_in == 8'hd2)? 32'h4410800e
	         : (byte_in == 8'hd3)? 32'h5af6029c
	         : (byte_in == 8'hd4)? 32'ha92d2a4b
	         : (byte_in == 8'hd5)? 32'hb7cba8d9
	         : (byte_in == 8'hd6)? 32'h79d9852a
	         : (byte_in == 8'hd7)? 32'h673f07b8
	         : (byte_in == 8'hd8)? 32'h350871ae
	         : (byte_in == 8'hd9)? 32'h2beef33c
	         : (byte_in == 8'hda)? 32'he5fcdecf
	         : (byte_in == 8'hdb)? 32'hfb1a5c5d
	         : (byte_in == 8'hdc)? 32'h08c1748a
	         : (byte_in == 8'hdd)? 32'h1627f618
	         : (byte_in == 8'hde)? 32'hd835dbeb
	         : (byte_in == 8'hdf)? 32'hc6d35979
	         : (byte_in == 8'he0)? 32'h4a93e323
	         : (byte_in == 8'he1)? 32'h547561b1
	         : (byte_in == 8'he2)? 32'h9a674c42
	         : (byte_in == 8'he3)? 32'h8481ced0
	         : (byte_in == 8'he4)? 32'h775ae607
	         : (byte_in == 8'he5)? 32'h69bc6495
	         : (byte_in == 8'he6)? 32'ha7ae4966
	         : (byte_in == 8'he7)? 32'hb948cbf4
	         : (byte_in == 8'he8)? 32'heb7fbde2
	         : (byte_in == 8'he9)? 32'hf5993f70
	         : (byte_in == 8'hea)? 32'h3b8b1283
	         : (byte_in == 8'heb)? 32'h256d9011
	         : (byte_in == 8'hec)? 32'hd6b6b8c6
	         : (byte_in == 8'hed)? 32'hc8503a54
	         : (byte_in == 8'hee)? 32'h064217a7
	         : (byte_in == 8'hef)? 32'h18a49535
	         : (byte_in == 8'hf0)? 32'h84a52f51
	         : (byte_in == 8'hf1)? 32'h9a43adc3
	         : (byte_in == 8'hf2)? 32'h54518030
	         : (byte_in == 8'hf3)? 32'h4ab702a2
	         : (byte_in == 8'hf4)? 32'hb96c2a75
	         : (byte_in == 8'hf5)? 32'ha78aa8e7
	         : (byte_in == 8'hf6)? 32'h69988514
	         : (byte_in == 8'hf7)? 32'h777e0786
	         : (byte_in == 8'hf8)? 32'h25497190
	         : (byte_in == 8'hf9)? 32'h3baff302
	         : (byte_in == 8'hfa)? 32'hf5bddef1
	         : (byte_in == 8'hfb)? 32'heb5b5c63
	         : (byte_in == 8'hfc)? 32'h188074b4
	         : (byte_in == 8'hfd)? 32'h0666f626
	         : (byte_in == 8'hfe)? 32'hc874dbd5
	         :                     32'hd6925947;

endmodule
//}}}

module TABLE16(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'hc8f10000
	         : (byte_in == 8'h02)? 32'h08bf0001
	         : (byte_in == 8'h03)? 32'hc04e0001
	         : (byte_in == 8'h04)? 32'h51ac0000
	         : (byte_in == 8'h05)? 32'h995d0000
	         : (byte_in == 8'h06)? 32'h59130001
	         : (byte_in == 8'h07)? 32'h91e20001
	         : (byte_in == 8'h08)? 32'hd98f0002
	         : (byte_in == 8'h09)? 32'h117e0002
	         : (byte_in == 8'h0a)? 32'hd1300003
	         : (byte_in == 8'h0b)? 32'h19c10003
	         : (byte_in == 8'h0c)? 32'h88230002
	         : (byte_in == 8'h0d)? 32'h40d20002
	         : (byte_in == 8'h0e)? 32'h809c0003
	         : (byte_in == 8'h0f)? 32'h486d0003
	         : (byte_in == 8'h10)? 32'h6ba90000
	         : (byte_in == 8'h11)? 32'ha3580000
	         : (byte_in == 8'h12)? 32'h63160001
	         : (byte_in == 8'h13)? 32'habe70001
	         : (byte_in == 8'h14)? 32'h3a050000
	         : (byte_in == 8'h15)? 32'hf2f40000
	         : (byte_in == 8'h16)? 32'h32ba0001
	         : (byte_in == 8'h17)? 32'hfa4b0001
	         : (byte_in == 8'h18)? 32'hb2260002
	         : (byte_in == 8'h19)? 32'h7ad70002
	         : (byte_in == 8'h1a)? 32'hba990003
	         : (byte_in == 8'h1b)? 32'h72680003
	         : (byte_in == 8'h1c)? 32'he38a0002
	         : (byte_in == 8'h1d)? 32'h2b7b0002
	         : (byte_in == 8'h1e)? 32'heb350003
	         : (byte_in == 8'h1f)? 32'h23c40003
	         : (byte_in == 8'h20)? 32'hbba10004
	         : (byte_in == 8'h21)? 32'h73500004
	         : (byte_in == 8'h22)? 32'hb31e0005
	         : (byte_in == 8'h23)? 32'h7bef0005
	         : (byte_in == 8'h24)? 32'hea0d0004
	         : (byte_in == 8'h25)? 32'h22fc0004
	         : (byte_in == 8'h26)? 32'he2b20005
	         : (byte_in == 8'h27)? 32'h2a430005
	         : (byte_in == 8'h28)? 32'h622e0006
	         : (byte_in == 8'h29)? 32'haadf0006
	         : (byte_in == 8'h2a)? 32'h6a910007
	         : (byte_in == 8'h2b)? 32'ha2600007
	         : (byte_in == 8'h2c)? 32'h33820006
	         : (byte_in == 8'h2d)? 32'hfb730006
	         : (byte_in == 8'h2e)? 32'h3b3d0007
	         : (byte_in == 8'h2f)? 32'hf3cc0007
	         : (byte_in == 8'h30)? 32'hd0080004
	         : (byte_in == 8'h31)? 32'h18f90004
	         : (byte_in == 8'h32)? 32'hd8b70005
	         : (byte_in == 8'h33)? 32'h10460005
	         : (byte_in == 8'h34)? 32'h81a40004
	         : (byte_in == 8'h35)? 32'h49550004
	         : (byte_in == 8'h36)? 32'h891b0005
	         : (byte_in == 8'h37)? 32'h41ea0005
	         : (byte_in == 8'h38)? 32'h09870006
	         : (byte_in == 8'h39)? 32'hc1760006
	         : (byte_in == 8'h3a)? 32'h01380007
	         : (byte_in == 8'h3b)? 32'hc9c90007
	         : (byte_in == 8'h3c)? 32'h582b0006
	         : (byte_in == 8'h3d)? 32'h90da0006
	         : (byte_in == 8'h3e)? 32'h50940007
	         : (byte_in == 8'h3f)? 32'h98650007
	         : (byte_in == 8'h40)? 32'h171c0000
	         : (byte_in == 8'h41)? 32'hdfed0000
	         : (byte_in == 8'h42)? 32'h1fa30001
	         : (byte_in == 8'h43)? 32'hd7520001
	         : (byte_in == 8'h44)? 32'h46b00000
	         : (byte_in == 8'h45)? 32'h8e410000
	         : (byte_in == 8'h46)? 32'h4e0f0001
	         : (byte_in == 8'h47)? 32'h86fe0001
	         : (byte_in == 8'h48)? 32'hce930002
	         : (byte_in == 8'h49)? 32'h06620002
	         : (byte_in == 8'h4a)? 32'hc62c0003
	         : (byte_in == 8'h4b)? 32'h0edd0003
	         : (byte_in == 8'h4c)? 32'h9f3f0002
	         : (byte_in == 8'h4d)? 32'h57ce0002
	         : (byte_in == 8'h4e)? 32'h97800003
	         : (byte_in == 8'h4f)? 32'h5f710003
	         : (byte_in == 8'h50)? 32'h7cb50000
	         : (byte_in == 8'h51)? 32'hb4440000
	         : (byte_in == 8'h52)? 32'h740a0001
	         : (byte_in == 8'h53)? 32'hbcfb0001
	         : (byte_in == 8'h54)? 32'h2d190000
	         : (byte_in == 8'h55)? 32'he5e80000
	         : (byte_in == 8'h56)? 32'h25a60001
	         : (byte_in == 8'h57)? 32'hed570001
	         : (byte_in == 8'h58)? 32'ha53a0002
	         : (byte_in == 8'h59)? 32'h6dcb0002
	         : (byte_in == 8'h5a)? 32'had850003
	         : (byte_in == 8'h5b)? 32'h65740003
	         : (byte_in == 8'h5c)? 32'hf4960002
	         : (byte_in == 8'h5d)? 32'h3c670002
	         : (byte_in == 8'h5e)? 32'hfc290003
	         : (byte_in == 8'h5f)? 32'h34d80003
	         : (byte_in == 8'h60)? 32'hacbd0004
	         : (byte_in == 8'h61)? 32'h644c0004
	         : (byte_in == 8'h62)? 32'ha4020005
	         : (byte_in == 8'h63)? 32'h6cf30005
	         : (byte_in == 8'h64)? 32'hfd110004
	         : (byte_in == 8'h65)? 32'h35e00004
	         : (byte_in == 8'h66)? 32'hf5ae0005
	         : (byte_in == 8'h67)? 32'h3d5f0005
	         : (byte_in == 8'h68)? 32'h75320006
	         : (byte_in == 8'h69)? 32'hbdc30006
	         : (byte_in == 8'h6a)? 32'h7d8d0007
	         : (byte_in == 8'h6b)? 32'hb57c0007
	         : (byte_in == 8'h6c)? 32'h249e0006
	         : (byte_in == 8'h6d)? 32'hec6f0006
	         : (byte_in == 8'h6e)? 32'h2c210007
	         : (byte_in == 8'h6f)? 32'he4d00007
	         : (byte_in == 8'h70)? 32'hc7140004
	         : (byte_in == 8'h71)? 32'h0fe50004
	         : (byte_in == 8'h72)? 32'hcfab0005
	         : (byte_in == 8'h73)? 32'h075a0005
	         : (byte_in == 8'h74)? 32'h96b80004
	         : (byte_in == 8'h75)? 32'h5e490004
	         : (byte_in == 8'h76)? 32'h9e070005
	         : (byte_in == 8'h77)? 32'h56f60005
	         : (byte_in == 8'h78)? 32'h1e9b0006
	         : (byte_in == 8'h79)? 32'hd66a0006
	         : (byte_in == 8'h7a)? 32'h16240007
	         : (byte_in == 8'h7b)? 32'hded50007
	         : (byte_in == 8'h7c)? 32'h4f370006
	         : (byte_in == 8'h7d)? 32'h87c60006
	         : (byte_in == 8'h7e)? 32'h47880007
	         : (byte_in == 8'h7f)? 32'h8f790007
	         : (byte_in == 8'h80)? 32'hbfb20008
	         : (byte_in == 8'h81)? 32'h77430008
	         : (byte_in == 8'h82)? 32'hb70d0009
	         : (byte_in == 8'h83)? 32'h7ffc0009
	         : (byte_in == 8'h84)? 32'hee1e0008
	         : (byte_in == 8'h85)? 32'h26ef0008
	         : (byte_in == 8'h86)? 32'he6a10009
	         : (byte_in == 8'h87)? 32'h2e500009
	         : (byte_in == 8'h88)? 32'h663d000a
	         : (byte_in == 8'h89)? 32'haecc000a
	         : (byte_in == 8'h8a)? 32'h6e82000b
	         : (byte_in == 8'h8b)? 32'ha673000b
	         : (byte_in == 8'h8c)? 32'h3791000a
	         : (byte_in == 8'h8d)? 32'hff60000a
	         : (byte_in == 8'h8e)? 32'h3f2e000b
	         : (byte_in == 8'h8f)? 32'hf7df000b
	         : (byte_in == 8'h90)? 32'hd41b0008
	         : (byte_in == 8'h91)? 32'h1cea0008
	         : (byte_in == 8'h92)? 32'hdca40009
	         : (byte_in == 8'h93)? 32'h14550009
	         : (byte_in == 8'h94)? 32'h85b70008
	         : (byte_in == 8'h95)? 32'h4d460008
	         : (byte_in == 8'h96)? 32'h8d080009
	         : (byte_in == 8'h97)? 32'h45f90009
	         : (byte_in == 8'h98)? 32'h0d94000a
	         : (byte_in == 8'h99)? 32'hc565000a
	         : (byte_in == 8'h9a)? 32'h052b000b
	         : (byte_in == 8'h9b)? 32'hcdda000b
	         : (byte_in == 8'h9c)? 32'h5c38000a
	         : (byte_in == 8'h9d)? 32'h94c9000a
	         : (byte_in == 8'h9e)? 32'h5487000b
	         : (byte_in == 8'h9f)? 32'h9c76000b
	         : (byte_in == 8'ha0)? 32'h0413000c
	         : (byte_in == 8'ha1)? 32'hcce2000c
	         : (byte_in == 8'ha2)? 32'h0cac000d
	         : (byte_in == 8'ha3)? 32'hc45d000d
	         : (byte_in == 8'ha4)? 32'h55bf000c
	         : (byte_in == 8'ha5)? 32'h9d4e000c
	         : (byte_in == 8'ha6)? 32'h5d00000d
	         : (byte_in == 8'ha7)? 32'h95f1000d
	         : (byte_in == 8'ha8)? 32'hdd9c000e
	         : (byte_in == 8'ha9)? 32'h156d000e
	         : (byte_in == 8'haa)? 32'hd523000f
	         : (byte_in == 8'hab)? 32'h1dd2000f
	         : (byte_in == 8'hac)? 32'h8c30000e
	         : (byte_in == 8'had)? 32'h44c1000e
	         : (byte_in == 8'hae)? 32'h848f000f
	         : (byte_in == 8'haf)? 32'h4c7e000f
	         : (byte_in == 8'hb0)? 32'h6fba000c
	         : (byte_in == 8'hb1)? 32'ha74b000c
	         : (byte_in == 8'hb2)? 32'h6705000d
	         : (byte_in == 8'hb3)? 32'haff4000d
	         : (byte_in == 8'hb4)? 32'h3e16000c
	         : (byte_in == 8'hb5)? 32'hf6e7000c
	         : (byte_in == 8'hb6)? 32'h36a9000d
	         : (byte_in == 8'hb7)? 32'hfe58000d
	         : (byte_in == 8'hb8)? 32'hb635000e
	         : (byte_in == 8'hb9)? 32'h7ec4000e
	         : (byte_in == 8'hba)? 32'hbe8a000f
	         : (byte_in == 8'hbb)? 32'h767b000f
	         : (byte_in == 8'hbc)? 32'he799000e
	         : (byte_in == 8'hbd)? 32'h2f68000e
	         : (byte_in == 8'hbe)? 32'hef26000f
	         : (byte_in == 8'hbf)? 32'h27d7000f
	         : (byte_in == 8'hc0)? 32'ha8ae0008
	         : (byte_in == 8'hc1)? 32'h605f0008
	         : (byte_in == 8'hc2)? 32'ha0110009
	         : (byte_in == 8'hc3)? 32'h68e00009
	         : (byte_in == 8'hc4)? 32'hf9020008
	         : (byte_in == 8'hc5)? 32'h31f30008
	         : (byte_in == 8'hc6)? 32'hf1bd0009
	         : (byte_in == 8'hc7)? 32'h394c0009
	         : (byte_in == 8'hc8)? 32'h7121000a
	         : (byte_in == 8'hc9)? 32'hb9d0000a
	         : (byte_in == 8'hca)? 32'h799e000b
	         : (byte_in == 8'hcb)? 32'hb16f000b
	         : (byte_in == 8'hcc)? 32'h208d000a
	         : (byte_in == 8'hcd)? 32'he87c000a
	         : (byte_in == 8'hce)? 32'h2832000b
	         : (byte_in == 8'hcf)? 32'he0c3000b
	         : (byte_in == 8'hd0)? 32'hc3070008
	         : (byte_in == 8'hd1)? 32'h0bf60008
	         : (byte_in == 8'hd2)? 32'hcbb80009
	         : (byte_in == 8'hd3)? 32'h03490009
	         : (byte_in == 8'hd4)? 32'h92ab0008
	         : (byte_in == 8'hd5)? 32'h5a5a0008
	         : (byte_in == 8'hd6)? 32'h9a140009
	         : (byte_in == 8'hd7)? 32'h52e50009
	         : (byte_in == 8'hd8)? 32'h1a88000a
	         : (byte_in == 8'hd9)? 32'hd279000a
	         : (byte_in == 8'hda)? 32'h1237000b
	         : (byte_in == 8'hdb)? 32'hdac6000b
	         : (byte_in == 8'hdc)? 32'h4b24000a
	         : (byte_in == 8'hdd)? 32'h83d5000a
	         : (byte_in == 8'hde)? 32'h439b000b
	         : (byte_in == 8'hdf)? 32'h8b6a000b
	         : (byte_in == 8'he0)? 32'h130f000c
	         : (byte_in == 8'he1)? 32'hdbfe000c
	         : (byte_in == 8'he2)? 32'h1bb0000d
	         : (byte_in == 8'he3)? 32'hd341000d
	         : (byte_in == 8'he4)? 32'h42a3000c
	         : (byte_in == 8'he5)? 32'h8a52000c
	         : (byte_in == 8'he6)? 32'h4a1c000d
	         : (byte_in == 8'he7)? 32'h82ed000d
	         : (byte_in == 8'he8)? 32'hca80000e
	         : (byte_in == 8'he9)? 32'h0271000e
	         : (byte_in == 8'hea)? 32'hc23f000f
	         : (byte_in == 8'heb)? 32'h0ace000f
	         : (byte_in == 8'hec)? 32'h9b2c000e
	         : (byte_in == 8'hed)? 32'h53dd000e
	         : (byte_in == 8'hee)? 32'h9393000f
	         : (byte_in == 8'hef)? 32'h5b62000f
	         : (byte_in == 8'hf0)? 32'h78a6000c
	         : (byte_in == 8'hf1)? 32'hb057000c
	         : (byte_in == 8'hf2)? 32'h7019000d
	         : (byte_in == 8'hf3)? 32'hb8e8000d
	         : (byte_in == 8'hf4)? 32'h290a000c
	         : (byte_in == 8'hf5)? 32'he1fb000c
	         : (byte_in == 8'hf6)? 32'h21b5000d
	         : (byte_in == 8'hf7)? 32'he944000d
	         : (byte_in == 8'hf8)? 32'ha129000e
	         : (byte_in == 8'hf9)? 32'h69d8000e
	         : (byte_in == 8'hfa)? 32'ha996000f
	         : (byte_in == 8'hfb)? 32'h6167000f
	         : (byte_in == 8'hfc)? 32'hf085000e
	         : (byte_in == 8'hfd)? 32'h3874000e
	         : (byte_in == 8'hfe)? 32'hf83a000f
	         :                     32'h30cb000f;

endmodule
//}}}

module TABLE17(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h2e390000
	         : (byte_in == 8'h02)? 32'h7f650010
	         : (byte_in == 8'h03)? 32'h515c0010
	         : (byte_in == 8'h04)? 32'h5c720000
	         : (byte_in == 8'h05)? 32'h724b0000
	         : (byte_in == 8'h06)? 32'h23170010
	         : (byte_in == 8'h07)? 32'h0d2e0010
	         : (byte_in == 8'h08)? 32'hfeca0020
	         : (byte_in == 8'h09)? 32'hd0f30020
	         : (byte_in == 8'h0a)? 32'h81af0030
	         : (byte_in == 8'h0b)? 32'haf960030
	         : (byte_in == 8'h0c)? 32'ha2b80020
	         : (byte_in == 8'h0d)? 32'h8c810020
	         : (byte_in == 8'h0e)? 32'hdddd0030
	         : (byte_in == 8'h0f)? 32'hf3e40030
	         : (byte_in == 8'h10)? 32'h78ab0000
	         : (byte_in == 8'h11)? 32'h56920000
	         : (byte_in == 8'h12)? 32'h07ce0010
	         : (byte_in == 8'h13)? 32'h29f70010
	         : (byte_in == 8'h14)? 32'h24d90000
	         : (byte_in == 8'h15)? 32'h0ae00000
	         : (byte_in == 8'h16)? 32'h5bbc0010
	         : (byte_in == 8'h17)? 32'h75850010
	         : (byte_in == 8'h18)? 32'h86610020
	         : (byte_in == 8'h19)? 32'ha8580020
	         : (byte_in == 8'h1a)? 32'hf9040030
	         : (byte_in == 8'h1b)? 32'hd73d0030
	         : (byte_in == 8'h1c)? 32'hda130020
	         : (byte_in == 8'h1d)? 32'hf42a0020
	         : (byte_in == 8'h1e)? 32'ha5760030
	         : (byte_in == 8'h1f)? 32'h8b4f0030
	         : (byte_in == 8'h20)? 32'h35650040
	         : (byte_in == 8'h21)? 32'h1b5c0040
	         : (byte_in == 8'h22)? 32'h4a000050
	         : (byte_in == 8'h23)? 32'h64390050
	         : (byte_in == 8'h24)? 32'h69170040
	         : (byte_in == 8'h25)? 32'h472e0040
	         : (byte_in == 8'h26)? 32'h16720050
	         : (byte_in == 8'h27)? 32'h384b0050
	         : (byte_in == 8'h28)? 32'hcbaf0060
	         : (byte_in == 8'h29)? 32'he5960060
	         : (byte_in == 8'h2a)? 32'hb4ca0070
	         : (byte_in == 8'h2b)? 32'h9af30070
	         : (byte_in == 8'h2c)? 32'h97dd0060
	         : (byte_in == 8'h2d)? 32'hb9e40060
	         : (byte_in == 8'h2e)? 32'he8b80070
	         : (byte_in == 8'h2f)? 32'hc6810070
	         : (byte_in == 8'h30)? 32'h4dce0040
	         : (byte_in == 8'h31)? 32'h63f70040
	         : (byte_in == 8'h32)? 32'h32ab0050
	         : (byte_in == 8'h33)? 32'h1c920050
	         : (byte_in == 8'h34)? 32'h11bc0040
	         : (byte_in == 8'h35)? 32'h3f850040
	         : (byte_in == 8'h36)? 32'h6ed90050
	         : (byte_in == 8'h37)? 32'h40e00050
	         : (byte_in == 8'h38)? 32'hb3040060
	         : (byte_in == 8'h39)? 32'h9d3d0060
	         : (byte_in == 8'h3a)? 32'hcc610070
	         : (byte_in == 8'h3b)? 32'he2580070
	         : (byte_in == 8'h3c)? 32'hef760060
	         : (byte_in == 8'h3d)? 32'hc14f0060
	         : (byte_in == 8'h3e)? 32'h90130070
	         : (byte_in == 8'h3f)? 32'hbe2a0070
	         : (byte_in == 8'h40)? 32'h39a60000
	         : (byte_in == 8'h41)? 32'h179f0000
	         : (byte_in == 8'h42)? 32'h46c30010
	         : (byte_in == 8'h43)? 32'h68fa0010
	         : (byte_in == 8'h44)? 32'h65d40000
	         : (byte_in == 8'h45)? 32'h4bed0000
	         : (byte_in == 8'h46)? 32'h1ab10010
	         : (byte_in == 8'h47)? 32'h34880010
	         : (byte_in == 8'h48)? 32'hc76c0020
	         : (byte_in == 8'h49)? 32'he9550020
	         : (byte_in == 8'h4a)? 32'hb8090030
	         : (byte_in == 8'h4b)? 32'h96300030
	         : (byte_in == 8'h4c)? 32'h9b1e0020
	         : (byte_in == 8'h4d)? 32'hb5270020
	         : (byte_in == 8'h4e)? 32'he47b0030
	         : (byte_in == 8'h4f)? 32'hca420030
	         : (byte_in == 8'h50)? 32'h410d0000
	         : (byte_in == 8'h51)? 32'h6f340000
	         : (byte_in == 8'h52)? 32'h3e680010
	         : (byte_in == 8'h53)? 32'h10510010
	         : (byte_in == 8'h54)? 32'h1d7f0000
	         : (byte_in == 8'h55)? 32'h33460000
	         : (byte_in == 8'h56)? 32'h621a0010
	         : (byte_in == 8'h57)? 32'h4c230010
	         : (byte_in == 8'h58)? 32'hbfc70020
	         : (byte_in == 8'h59)? 32'h91fe0020
	         : (byte_in == 8'h5a)? 32'hc0a20030
	         : (byte_in == 8'h5b)? 32'hee9b0030
	         : (byte_in == 8'h5c)? 32'he3b50020
	         : (byte_in == 8'h5d)? 32'hcd8c0020
	         : (byte_in == 8'h5e)? 32'h9cd00030
	         : (byte_in == 8'h5f)? 32'hb2e90030
	         : (byte_in == 8'h60)? 32'h0cc30040
	         : (byte_in == 8'h61)? 32'h22fa0040
	         : (byte_in == 8'h62)? 32'h73a60050
	         : (byte_in == 8'h63)? 32'h5d9f0050
	         : (byte_in == 8'h64)? 32'h50b10040
	         : (byte_in == 8'h65)? 32'h7e880040
	         : (byte_in == 8'h66)? 32'h2fd40050
	         : (byte_in == 8'h67)? 32'h01ed0050
	         : (byte_in == 8'h68)? 32'hf2090060
	         : (byte_in == 8'h69)? 32'hdc300060
	         : (byte_in == 8'h6a)? 32'h8d6c0070
	         : (byte_in == 8'h6b)? 32'ha3550070
	         : (byte_in == 8'h6c)? 32'hae7b0060
	         : (byte_in == 8'h6d)? 32'h80420060
	         : (byte_in == 8'h6e)? 32'hd11e0070
	         : (byte_in == 8'h6f)? 32'hff270070
	         : (byte_in == 8'h70)? 32'h74680040
	         : (byte_in == 8'h71)? 32'h5a510040
	         : (byte_in == 8'h72)? 32'h0b0d0050
	         : (byte_in == 8'h73)? 32'h25340050
	         : (byte_in == 8'h74)? 32'h281a0040
	         : (byte_in == 8'h75)? 32'h06230040
	         : (byte_in == 8'h76)? 32'h577f0050
	         : (byte_in == 8'h77)? 32'h79460050
	         : (byte_in == 8'h78)? 32'h8aa20060
	         : (byte_in == 8'h79)? 32'ha49b0060
	         : (byte_in == 8'h7a)? 32'hf5c70070
	         : (byte_in == 8'h7b)? 32'hdbfe0070
	         : (byte_in == 8'h7c)? 32'hd6d00060
	         : (byte_in == 8'h7d)? 32'hf8e90060
	         : (byte_in == 8'h7e)? 32'ha9b50070
	         : (byte_in == 8'h7f)? 32'h878c0070
	         : (byte_in == 8'h80)? 32'h62740080
	         : (byte_in == 8'h81)? 32'h4c4d0080
	         : (byte_in == 8'h82)? 32'h1d110090
	         : (byte_in == 8'h83)? 32'h33280090
	         : (byte_in == 8'h84)? 32'h3e060080
	         : (byte_in == 8'h85)? 32'h103f0080
	         : (byte_in == 8'h86)? 32'h41630090
	         : (byte_in == 8'h87)? 32'h6f5a0090
	         : (byte_in == 8'h88)? 32'h9cbe00a0
	         : (byte_in == 8'h89)? 32'hb28700a0
	         : (byte_in == 8'h8a)? 32'he3db00b0
	         : (byte_in == 8'h8b)? 32'hcde200b0
	         : (byte_in == 8'h8c)? 32'hc0cc00a0
	         : (byte_in == 8'h8d)? 32'heef500a0
	         : (byte_in == 8'h8e)? 32'hbfa900b0
	         : (byte_in == 8'h8f)? 32'h919000b0
	         : (byte_in == 8'h90)? 32'h1adf0080
	         : (byte_in == 8'h91)? 32'h34e60080
	         : (byte_in == 8'h92)? 32'h65ba0090
	         : (byte_in == 8'h93)? 32'h4b830090
	         : (byte_in == 8'h94)? 32'h46ad0080
	         : (byte_in == 8'h95)? 32'h68940080
	         : (byte_in == 8'h96)? 32'h39c80090
	         : (byte_in == 8'h97)? 32'h17f10090
	         : (byte_in == 8'h98)? 32'he41500a0
	         : (byte_in == 8'h99)? 32'hca2c00a0
	         : (byte_in == 8'h9a)? 32'h9b7000b0
	         : (byte_in == 8'h9b)? 32'hb54900b0
	         : (byte_in == 8'h9c)? 32'hb86700a0
	         : (byte_in == 8'h9d)? 32'h965e00a0
	         : (byte_in == 8'h9e)? 32'hc70200b0
	         : (byte_in == 8'h9f)? 32'he93b00b0
	         : (byte_in == 8'ha0)? 32'h571100c0
	         : (byte_in == 8'ha1)? 32'h792800c0
	         : (byte_in == 8'ha2)? 32'h287400d0
	         : (byte_in == 8'ha3)? 32'h064d00d0
	         : (byte_in == 8'ha4)? 32'h0b6300c0
	         : (byte_in == 8'ha5)? 32'h255a00c0
	         : (byte_in == 8'ha6)? 32'h740600d0
	         : (byte_in == 8'ha7)? 32'h5a3f00d0
	         : (byte_in == 8'ha8)? 32'ha9db00e0
	         : (byte_in == 8'ha9)? 32'h87e200e0
	         : (byte_in == 8'haa)? 32'hd6be00f0
	         : (byte_in == 8'hab)? 32'hf88700f0
	         : (byte_in == 8'hac)? 32'hf5a900e0
	         : (byte_in == 8'had)? 32'hdb9000e0
	         : (byte_in == 8'hae)? 32'h8acc00f0
	         : (byte_in == 8'haf)? 32'ha4f500f0
	         : (byte_in == 8'hb0)? 32'h2fba00c0
	         : (byte_in == 8'hb1)? 32'h018300c0
	         : (byte_in == 8'hb2)? 32'h50df00d0
	         : (byte_in == 8'hb3)? 32'h7ee600d0
	         : (byte_in == 8'hb4)? 32'h73c800c0
	         : (byte_in == 8'hb5)? 32'h5df100c0
	         : (byte_in == 8'hb6)? 32'h0cad00d0
	         : (byte_in == 8'hb7)? 32'h229400d0
	         : (byte_in == 8'hb8)? 32'hd17000e0
	         : (byte_in == 8'hb9)? 32'hff4900e0
	         : (byte_in == 8'hba)? 32'hae1500f0
	         : (byte_in == 8'hbb)? 32'h802c00f0
	         : (byte_in == 8'hbc)? 32'h8d0200e0
	         : (byte_in == 8'hbd)? 32'ha33b00e0
	         : (byte_in == 8'hbe)? 32'hf26700f0
	         : (byte_in == 8'hbf)? 32'hdc5e00f0
	         : (byte_in == 8'hc0)? 32'h5bd20080
	         : (byte_in == 8'hc1)? 32'h75eb0080
	         : (byte_in == 8'hc2)? 32'h24b70090
	         : (byte_in == 8'hc3)? 32'h0a8e0090
	         : (byte_in == 8'hc4)? 32'h07a00080
	         : (byte_in == 8'hc5)? 32'h29990080
	         : (byte_in == 8'hc6)? 32'h78c50090
	         : (byte_in == 8'hc7)? 32'h56fc0090
	         : (byte_in == 8'hc8)? 32'ha51800a0
	         : (byte_in == 8'hc9)? 32'h8b2100a0
	         : (byte_in == 8'hca)? 32'hda7d00b0
	         : (byte_in == 8'hcb)? 32'hf44400b0
	         : (byte_in == 8'hcc)? 32'hf96a00a0
	         : (byte_in == 8'hcd)? 32'hd75300a0
	         : (byte_in == 8'hce)? 32'h860f00b0
	         : (byte_in == 8'hcf)? 32'ha83600b0
	         : (byte_in == 8'hd0)? 32'h23790080
	         : (byte_in == 8'hd1)? 32'h0d400080
	         : (byte_in == 8'hd2)? 32'h5c1c0090
	         : (byte_in == 8'hd3)? 32'h72250090
	         : (byte_in == 8'hd4)? 32'h7f0b0080
	         : (byte_in == 8'hd5)? 32'h51320080
	         : (byte_in == 8'hd6)? 32'h006e0090
	         : (byte_in == 8'hd7)? 32'h2e570090
	         : (byte_in == 8'hd8)? 32'hddb300a0
	         : (byte_in == 8'hd9)? 32'hf38a00a0
	         : (byte_in == 8'hda)? 32'ha2d600b0
	         : (byte_in == 8'hdb)? 32'h8cef00b0
	         : (byte_in == 8'hdc)? 32'h81c100a0
	         : (byte_in == 8'hdd)? 32'haff800a0
	         : (byte_in == 8'hde)? 32'hfea400b0
	         : (byte_in == 8'hdf)? 32'hd09d00b0
	         : (byte_in == 8'he0)? 32'h6eb700c0
	         : (byte_in == 8'he1)? 32'h408e00c0
	         : (byte_in == 8'he2)? 32'h11d200d0
	         : (byte_in == 8'he3)? 32'h3feb00d0
	         : (byte_in == 8'he4)? 32'h32c500c0
	         : (byte_in == 8'he5)? 32'h1cfc00c0
	         : (byte_in == 8'he6)? 32'h4da000d0
	         : (byte_in == 8'he7)? 32'h639900d0
	         : (byte_in == 8'he8)? 32'h907d00e0
	         : (byte_in == 8'he9)? 32'hbe4400e0
	         : (byte_in == 8'hea)? 32'hef1800f0
	         : (byte_in == 8'heb)? 32'hc12100f0
	         : (byte_in == 8'hec)? 32'hcc0f00e0
	         : (byte_in == 8'hed)? 32'he23600e0
	         : (byte_in == 8'hee)? 32'hb36a00f0
	         : (byte_in == 8'hef)? 32'h9d5300f0
	         : (byte_in == 8'hf0)? 32'h161c00c0
	         : (byte_in == 8'hf1)? 32'h382500c0
	         : (byte_in == 8'hf2)? 32'h697900d0
	         : (byte_in == 8'hf3)? 32'h474000d0
	         : (byte_in == 8'hf4)? 32'h4a6e00c0
	         : (byte_in == 8'hf5)? 32'h645700c0
	         : (byte_in == 8'hf6)? 32'h350b00d0
	         : (byte_in == 8'hf7)? 32'h1b3200d0
	         : (byte_in == 8'hf8)? 32'he8d600e0
	         : (byte_in == 8'hf9)? 32'hc6ef00e0
	         : (byte_in == 8'hfa)? 32'h97b300f0
	         : (byte_in == 8'hfb)? 32'hb98a00f0
	         : (byte_in == 8'hfc)? 32'hb4a400e0
	         : (byte_in == 8'hfd)? 32'h9a9d00e0
	         : (byte_in == 8'hfe)? 32'hcbc100f0
	         :                     32'he5f800f0;

endmodule
//}}}

module TABLE18(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h734c0000
	         : (byte_in == 8'h02)? 32'hc4e80100
	         : (byte_in == 8'h03)? 32'hb7a40100
	         : (byte_in == 8'h04)? 32'hee260000
	         : (byte_in == 8'h05)? 32'h9d6a0000
	         : (byte_in == 8'h06)? 32'h2ace0100
	         : (byte_in == 8'h07)? 32'h59820100
	         : (byte_in == 8'h08)? 32'h499e0200
	         : (byte_in == 8'h09)? 32'h3ad20200
	         : (byte_in == 8'h0a)? 32'h8d760300
	         : (byte_in == 8'h0b)? 32'hfe3a0300
	         : (byte_in == 8'h0c)? 32'ha7b80200
	         : (byte_in == 8'h0d)? 32'hd4f40200
	         : (byte_in == 8'h0e)? 32'h63500300
	         : (byte_in == 8'h0f)? 32'h101c0300
	         : (byte_in == 8'h10)? 32'h14bd0000
	         : (byte_in == 8'h11)? 32'h67f10000
	         : (byte_in == 8'h12)? 32'hd0550100
	         : (byte_in == 8'h13)? 32'ha3190100
	         : (byte_in == 8'h14)? 32'hfa9b0000
	         : (byte_in == 8'h15)? 32'h89d70000
	         : (byte_in == 8'h16)? 32'h3e730100
	         : (byte_in == 8'h17)? 32'h4d3f0100
	         : (byte_in == 8'h18)? 32'h5d230200
	         : (byte_in == 8'h19)? 32'h2e6f0200
	         : (byte_in == 8'h1a)? 32'h99cb0300
	         : (byte_in == 8'h1b)? 32'hea870300
	         : (byte_in == 8'h1c)? 32'hb3050200
	         : (byte_in == 8'h1d)? 32'hc0490200
	         : (byte_in == 8'h1e)? 32'h77ed0300
	         : (byte_in == 8'h1f)? 32'h04a10300
	         : (byte_in == 8'h20)? 32'h9b830400
	         : (byte_in == 8'h21)? 32'he8cf0400
	         : (byte_in == 8'h22)? 32'h5f6b0500
	         : (byte_in == 8'h23)? 32'h2c270500
	         : (byte_in == 8'h24)? 32'h75a50400
	         : (byte_in == 8'h25)? 32'h06e90400
	         : (byte_in == 8'h26)? 32'hb14d0500
	         : (byte_in == 8'h27)? 32'hc2010500
	         : (byte_in == 8'h28)? 32'hd21d0600
	         : (byte_in == 8'h29)? 32'ha1510600
	         : (byte_in == 8'h2a)? 32'h16f50700
	         : (byte_in == 8'h2b)? 32'h65b90700
	         : (byte_in == 8'h2c)? 32'h3c3b0600
	         : (byte_in == 8'h2d)? 32'h4f770600
	         : (byte_in == 8'h2e)? 32'hf8d30700
	         : (byte_in == 8'h2f)? 32'h8b9f0700
	         : (byte_in == 8'h30)? 32'h8f3e0400
	         : (byte_in == 8'h31)? 32'hfc720400
	         : (byte_in == 8'h32)? 32'h4bd60500
	         : (byte_in == 8'h33)? 32'h389a0500
	         : (byte_in == 8'h34)? 32'h61180400
	         : (byte_in == 8'h35)? 32'h12540400
	         : (byte_in == 8'h36)? 32'ha5f00500
	         : (byte_in == 8'h37)? 32'hd6bc0500
	         : (byte_in == 8'h38)? 32'hc6a00600
	         : (byte_in == 8'h39)? 32'hb5ec0600
	         : (byte_in == 8'h3a)? 32'h02480700
	         : (byte_in == 8'h3b)? 32'h71040700
	         : (byte_in == 8'h3c)? 32'h28860600
	         : (byte_in == 8'h3d)? 32'h5bca0600
	         : (byte_in == 8'h3e)? 32'hec6e0700
	         : (byte_in == 8'h3f)? 32'h9f220700
	         : (byte_in == 8'h40)? 32'he18b0000
	         : (byte_in == 8'h41)? 32'h92c70000
	         : (byte_in == 8'h42)? 32'h25630100
	         : (byte_in == 8'h43)? 32'h562f0100
	         : (byte_in == 8'h44)? 32'h0fad0000
	         : (byte_in == 8'h45)? 32'h7ce10000
	         : (byte_in == 8'h46)? 32'hcb450100
	         : (byte_in == 8'h47)? 32'hb8090100
	         : (byte_in == 8'h48)? 32'ha8150200
	         : (byte_in == 8'h49)? 32'hdb590200
	         : (byte_in == 8'h4a)? 32'h6cfd0300
	         : (byte_in == 8'h4b)? 32'h1fb10300
	         : (byte_in == 8'h4c)? 32'h46330200
	         : (byte_in == 8'h4d)? 32'h357f0200
	         : (byte_in == 8'h4e)? 32'h82db0300
	         : (byte_in == 8'h4f)? 32'hf1970300
	         : (byte_in == 8'h50)? 32'hf5360000
	         : (byte_in == 8'h51)? 32'h867a0000
	         : (byte_in == 8'h52)? 32'h31de0100
	         : (byte_in == 8'h53)? 32'h42920100
	         : (byte_in == 8'h54)? 32'h1b100000
	         : (byte_in == 8'h55)? 32'h685c0000
	         : (byte_in == 8'h56)? 32'hdff80100
	         : (byte_in == 8'h57)? 32'hacb40100
	         : (byte_in == 8'h58)? 32'hbca80200
	         : (byte_in == 8'h59)? 32'hcfe40200
	         : (byte_in == 8'h5a)? 32'h78400300
	         : (byte_in == 8'h5b)? 32'h0b0c0300
	         : (byte_in == 8'h5c)? 32'h528e0200
	         : (byte_in == 8'h5d)? 32'h21c20200
	         : (byte_in == 8'h5e)? 32'h96660300
	         : (byte_in == 8'h5f)? 32'he52a0300
	         : (byte_in == 8'h60)? 32'h7a080400
	         : (byte_in == 8'h61)? 32'h09440400
	         : (byte_in == 8'h62)? 32'hbee00500
	         : (byte_in == 8'h63)? 32'hcdac0500
	         : (byte_in == 8'h64)? 32'h942e0400
	         : (byte_in == 8'h65)? 32'he7620400
	         : (byte_in == 8'h66)? 32'h50c60500
	         : (byte_in == 8'h67)? 32'h238a0500
	         : (byte_in == 8'h68)? 32'h33960600
	         : (byte_in == 8'h69)? 32'h40da0600
	         : (byte_in == 8'h6a)? 32'hf77e0700
	         : (byte_in == 8'h6b)? 32'h84320700
	         : (byte_in == 8'h6c)? 32'hddb00600
	         : (byte_in == 8'h6d)? 32'haefc0600
	         : (byte_in == 8'h6e)? 32'h19580700
	         : (byte_in == 8'h6f)? 32'h6a140700
	         : (byte_in == 8'h70)? 32'h6eb50400
	         : (byte_in == 8'h71)? 32'h1df90400
	         : (byte_in == 8'h72)? 32'haa5d0500
	         : (byte_in == 8'h73)? 32'hd9110500
	         : (byte_in == 8'h74)? 32'h80930400
	         : (byte_in == 8'h75)? 32'hf3df0400
	         : (byte_in == 8'h76)? 32'h447b0500
	         : (byte_in == 8'h77)? 32'h37370500
	         : (byte_in == 8'h78)? 32'h272b0600
	         : (byte_in == 8'h79)? 32'h54670600
	         : (byte_in == 8'h7a)? 32'he3c30700
	         : (byte_in == 8'h7b)? 32'h908f0700
	         : (byte_in == 8'h7c)? 32'hc90d0600
	         : (byte_in == 8'h7d)? 32'hba410600
	         : (byte_in == 8'h7e)? 32'h0de50700
	         : (byte_in == 8'h7f)? 32'h7ea90700
	         : (byte_in == 8'h80)? 32'h3fb90800
	         : (byte_in == 8'h81)? 32'h4cf50800
	         : (byte_in == 8'h82)? 32'hfb510900
	         : (byte_in == 8'h83)? 32'h881d0900
	         : (byte_in == 8'h84)? 32'hd19f0800
	         : (byte_in == 8'h85)? 32'ha2d30800
	         : (byte_in == 8'h86)? 32'h15770900
	         : (byte_in == 8'h87)? 32'h663b0900
	         : (byte_in == 8'h88)? 32'h76270a00
	         : (byte_in == 8'h89)? 32'h056b0a00
	         : (byte_in == 8'h8a)? 32'hb2cf0b00
	         : (byte_in == 8'h8b)? 32'hc1830b00
	         : (byte_in == 8'h8c)? 32'h98010a00
	         : (byte_in == 8'h8d)? 32'heb4d0a00
	         : (byte_in == 8'h8e)? 32'h5ce90b00
	         : (byte_in == 8'h8f)? 32'h2fa50b00
	         : (byte_in == 8'h90)? 32'h2b040800
	         : (byte_in == 8'h91)? 32'h58480800
	         : (byte_in == 8'h92)? 32'hefec0900
	         : (byte_in == 8'h93)? 32'h9ca00900
	         : (byte_in == 8'h94)? 32'hc5220800
	         : (byte_in == 8'h95)? 32'hb66e0800
	         : (byte_in == 8'h96)? 32'h01ca0900
	         : (byte_in == 8'h97)? 32'h72860900
	         : (byte_in == 8'h98)? 32'h629a0a00
	         : (byte_in == 8'h99)? 32'h11d60a00
	         : (byte_in == 8'h9a)? 32'ha6720b00
	         : (byte_in == 8'h9b)? 32'hd53e0b00
	         : (byte_in == 8'h9c)? 32'h8cbc0a00
	         : (byte_in == 8'h9d)? 32'hfff00a00
	         : (byte_in == 8'h9e)? 32'h48540b00
	         : (byte_in == 8'h9f)? 32'h3b180b00
	         : (byte_in == 8'ha0)? 32'ha43a0c00
	         : (byte_in == 8'ha1)? 32'hd7760c00
	         : (byte_in == 8'ha2)? 32'h60d20d00
	         : (byte_in == 8'ha3)? 32'h139e0d00
	         : (byte_in == 8'ha4)? 32'h4a1c0c00
	         : (byte_in == 8'ha5)? 32'h39500c00
	         : (byte_in == 8'ha6)? 32'h8ef40d00
	         : (byte_in == 8'ha7)? 32'hfdb80d00
	         : (byte_in == 8'ha8)? 32'heda40e00
	         : (byte_in == 8'ha9)? 32'h9ee80e00
	         : (byte_in == 8'haa)? 32'h294c0f00
	         : (byte_in == 8'hab)? 32'h5a000f00
	         : (byte_in == 8'hac)? 32'h03820e00
	         : (byte_in == 8'had)? 32'h70ce0e00
	         : (byte_in == 8'hae)? 32'hc76a0f00
	         : (byte_in == 8'haf)? 32'hb4260f00
	         : (byte_in == 8'hb0)? 32'hb0870c00
	         : (byte_in == 8'hb1)? 32'hc3cb0c00
	         : (byte_in == 8'hb2)? 32'h746f0d00
	         : (byte_in == 8'hb3)? 32'h07230d00
	         : (byte_in == 8'hb4)? 32'h5ea10c00
	         : (byte_in == 8'hb5)? 32'h2ded0c00
	         : (byte_in == 8'hb6)? 32'h9a490d00
	         : (byte_in == 8'hb7)? 32'he9050d00
	         : (byte_in == 8'hb8)? 32'hf9190e00
	         : (byte_in == 8'hb9)? 32'h8a550e00
	         : (byte_in == 8'hba)? 32'h3df10f00
	         : (byte_in == 8'hbb)? 32'h4ebd0f00
	         : (byte_in == 8'hbc)? 32'h173f0e00
	         : (byte_in == 8'hbd)? 32'h64730e00
	         : (byte_in == 8'hbe)? 32'hd3d70f00
	         : (byte_in == 8'hbf)? 32'ha09b0f00
	         : (byte_in == 8'hc0)? 32'hde320800
	         : (byte_in == 8'hc1)? 32'had7e0800
	         : (byte_in == 8'hc2)? 32'h1ada0900
	         : (byte_in == 8'hc3)? 32'h69960900
	         : (byte_in == 8'hc4)? 32'h30140800
	         : (byte_in == 8'hc5)? 32'h43580800
	         : (byte_in == 8'hc6)? 32'hf4fc0900
	         : (byte_in == 8'hc7)? 32'h87b00900
	         : (byte_in == 8'hc8)? 32'h97ac0a00
	         : (byte_in == 8'hc9)? 32'he4e00a00
	         : (byte_in == 8'hca)? 32'h53440b00
	         : (byte_in == 8'hcb)? 32'h20080b00
	         : (byte_in == 8'hcc)? 32'h798a0a00
	         : (byte_in == 8'hcd)? 32'h0ac60a00
	         : (byte_in == 8'hce)? 32'hbd620b00
	         : (byte_in == 8'hcf)? 32'hce2e0b00
	         : (byte_in == 8'hd0)? 32'hca8f0800
	         : (byte_in == 8'hd1)? 32'hb9c30800
	         : (byte_in == 8'hd2)? 32'h0e670900
	         : (byte_in == 8'hd3)? 32'h7d2b0900
	         : (byte_in == 8'hd4)? 32'h24a90800
	         : (byte_in == 8'hd5)? 32'h57e50800
	         : (byte_in == 8'hd6)? 32'he0410900
	         : (byte_in == 8'hd7)? 32'h930d0900
	         : (byte_in == 8'hd8)? 32'h83110a00
	         : (byte_in == 8'hd9)? 32'hf05d0a00
	         : (byte_in == 8'hda)? 32'h47f90b00
	         : (byte_in == 8'hdb)? 32'h34b50b00
	         : (byte_in == 8'hdc)? 32'h6d370a00
	         : (byte_in == 8'hdd)? 32'h1e7b0a00
	         : (byte_in == 8'hde)? 32'ha9df0b00
	         : (byte_in == 8'hdf)? 32'hda930b00
	         : (byte_in == 8'he0)? 32'h45b10c00
	         : (byte_in == 8'he1)? 32'h36fd0c00
	         : (byte_in == 8'he2)? 32'h81590d00
	         : (byte_in == 8'he3)? 32'hf2150d00
	         : (byte_in == 8'he4)? 32'hab970c00
	         : (byte_in == 8'he5)? 32'hd8db0c00
	         : (byte_in == 8'he6)? 32'h6f7f0d00
	         : (byte_in == 8'he7)? 32'h1c330d00
	         : (byte_in == 8'he8)? 32'h0c2f0e00
	         : (byte_in == 8'he9)? 32'h7f630e00
	         : (byte_in == 8'hea)? 32'hc8c70f00
	         : (byte_in == 8'heb)? 32'hbb8b0f00
	         : (byte_in == 8'hec)? 32'he2090e00
	         : (byte_in == 8'hed)? 32'h91450e00
	         : (byte_in == 8'hee)? 32'h26e10f00
	         : (byte_in == 8'hef)? 32'h55ad0f00
	         : (byte_in == 8'hf0)? 32'h510c0c00
	         : (byte_in == 8'hf1)? 32'h22400c00
	         : (byte_in == 8'hf2)? 32'h95e40d00
	         : (byte_in == 8'hf3)? 32'he6a80d00
	         : (byte_in == 8'hf4)? 32'hbf2a0c00
	         : (byte_in == 8'hf5)? 32'hcc660c00
	         : (byte_in == 8'hf6)? 32'h7bc20d00
	         : (byte_in == 8'hf7)? 32'h088e0d00
	         : (byte_in == 8'hf8)? 32'h18920e00
	         : (byte_in == 8'hf9)? 32'h6bde0e00
	         : (byte_in == 8'hfa)? 32'hdc7a0f00
	         : (byte_in == 8'hfb)? 32'haf360f00
	         : (byte_in == 8'hfc)? 32'hf6b40e00
	         : (byte_in == 8'hfd)? 32'h85f80e00
	         : (byte_in == 8'hfe)? 32'h325c0f00
	         :                     32'h41100f00;

endmodule
//}}}

module TABLE19(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'hcba90000
	         : (byte_in == 8'h02)? 32'hbf3c1000
	         : (byte_in == 8'h03)? 32'h74951000
	         : (byte_in == 8'h04)? 32'h97530000
	         : (byte_in == 8'h05)? 32'h5cfa0000
	         : (byte_in == 8'h06)? 32'h286f1000
	         : (byte_in == 8'h07)? 32'he3c61000
	         : (byte_in == 8'h08)? 32'h7e792000
	         : (byte_in == 8'h09)? 32'hb5d02000
	         : (byte_in == 8'h0a)? 32'hc1453000
	         : (byte_in == 8'h0b)? 32'h0aec3000
	         : (byte_in == 8'h0c)? 32'he92a2000
	         : (byte_in == 8'h0d)? 32'h22832000
	         : (byte_in == 8'h0e)? 32'h56163000
	         : (byte_in == 8'h0f)? 32'h9dbf3000
	         : (byte_in == 8'h10)? 32'he6570000
	         : (byte_in == 8'h11)? 32'h2dfe0000
	         : (byte_in == 8'h12)? 32'h596b1000
	         : (byte_in == 8'h13)? 32'h92c21000
	         : (byte_in == 8'h14)? 32'h71040000
	         : (byte_in == 8'h15)? 32'hbaad0000
	         : (byte_in == 8'h16)? 32'hce381000
	         : (byte_in == 8'h17)? 32'h05911000
	         : (byte_in == 8'h18)? 32'h982e2000
	         : (byte_in == 8'h19)? 32'h53872000
	         : (byte_in == 8'h1a)? 32'h27123000
	         : (byte_in == 8'h1b)? 32'hecbb3000
	         : (byte_in == 8'h1c)? 32'h0f7d2000
	         : (byte_in == 8'h1d)? 32'hc4d42000
	         : (byte_in == 8'h1e)? 32'hb0413000
	         : (byte_in == 8'h1f)? 32'h7be83000
	         : (byte_in == 8'h20)? 32'hf44c4000
	         : (byte_in == 8'h21)? 32'h3fe54000
	         : (byte_in == 8'h22)? 32'h4b705000
	         : (byte_in == 8'h23)? 32'h80d95000
	         : (byte_in == 8'h24)? 32'h631f4000
	         : (byte_in == 8'h25)? 32'ha8b64000
	         : (byte_in == 8'h26)? 32'hdc235000
	         : (byte_in == 8'h27)? 32'h178a5000
	         : (byte_in == 8'h28)? 32'h8a356000
	         : (byte_in == 8'h29)? 32'h419c6000
	         : (byte_in == 8'h2a)? 32'h35097000
	         : (byte_in == 8'h2b)? 32'hfea07000
	         : (byte_in == 8'h2c)? 32'h1d666000
	         : (byte_in == 8'h2d)? 32'hd6cf6000
	         : (byte_in == 8'h2e)? 32'ha25a7000
	         : (byte_in == 8'h2f)? 32'h69f37000
	         : (byte_in == 8'h30)? 32'h121b4000
	         : (byte_in == 8'h31)? 32'hd9b24000
	         : (byte_in == 8'h32)? 32'had275000
	         : (byte_in == 8'h33)? 32'h668e5000
	         : (byte_in == 8'h34)? 32'h85484000
	         : (byte_in == 8'h35)? 32'h4ee14000
	         : (byte_in == 8'h36)? 32'h3a745000
	         : (byte_in == 8'h37)? 32'hf1dd5000
	         : (byte_in == 8'h38)? 32'h6c626000
	         : (byte_in == 8'h39)? 32'ha7cb6000
	         : (byte_in == 8'h3a)? 32'hd35e7000
	         : (byte_in == 8'h3b)? 32'h18f77000
	         : (byte_in == 8'h3c)? 32'hfb316000
	         : (byte_in == 8'h3d)? 32'h30986000
	         : (byte_in == 8'h3e)? 32'h440d7000
	         : (byte_in == 8'h3f)? 32'h8fa47000
	         : (byte_in == 8'h40)? 32'h045f0000
	         : (byte_in == 8'h41)? 32'hcff60000
	         : (byte_in == 8'h42)? 32'hbb631000
	         : (byte_in == 8'h43)? 32'h70ca1000
	         : (byte_in == 8'h44)? 32'h930c0000
	         : (byte_in == 8'h45)? 32'h58a50000
	         : (byte_in == 8'h46)? 32'h2c301000
	         : (byte_in == 8'h47)? 32'he7991000
	         : (byte_in == 8'h48)? 32'h7a262000
	         : (byte_in == 8'h49)? 32'hb18f2000
	         : (byte_in == 8'h4a)? 32'hc51a3000
	         : (byte_in == 8'h4b)? 32'h0eb33000
	         : (byte_in == 8'h4c)? 32'hed752000
	         : (byte_in == 8'h4d)? 32'h26dc2000
	         : (byte_in == 8'h4e)? 32'h52493000
	         : (byte_in == 8'h4f)? 32'h99e03000
	         : (byte_in == 8'h50)? 32'he2080000
	         : (byte_in == 8'h51)? 32'h29a10000
	         : (byte_in == 8'h52)? 32'h5d341000
	         : (byte_in == 8'h53)? 32'h969d1000
	         : (byte_in == 8'h54)? 32'h755b0000
	         : (byte_in == 8'h55)? 32'hbef20000
	         : (byte_in == 8'h56)? 32'hca671000
	         : (byte_in == 8'h57)? 32'h01ce1000
	         : (byte_in == 8'h58)? 32'h9c712000
	         : (byte_in == 8'h59)? 32'h57d82000
	         : (byte_in == 8'h5a)? 32'h234d3000
	         : (byte_in == 8'h5b)? 32'he8e43000
	         : (byte_in == 8'h5c)? 32'h0b222000
	         : (byte_in == 8'h5d)? 32'hc08b2000
	         : (byte_in == 8'h5e)? 32'hb41e3000
	         : (byte_in == 8'h5f)? 32'h7fb73000
	         : (byte_in == 8'h60)? 32'hf0134000
	         : (byte_in == 8'h61)? 32'h3bba4000
	         : (byte_in == 8'h62)? 32'h4f2f5000
	         : (byte_in == 8'h63)? 32'h84865000
	         : (byte_in == 8'h64)? 32'h67404000
	         : (byte_in == 8'h65)? 32'hace94000
	         : (byte_in == 8'h66)? 32'hd87c5000
	         : (byte_in == 8'h67)? 32'h13d55000
	         : (byte_in == 8'h68)? 32'h8e6a6000
	         : (byte_in == 8'h69)? 32'h45c36000
	         : (byte_in == 8'h6a)? 32'h31567000
	         : (byte_in == 8'h6b)? 32'hfaff7000
	         : (byte_in == 8'h6c)? 32'h19396000
	         : (byte_in == 8'h6d)? 32'hd2906000
	         : (byte_in == 8'h6e)? 32'ha6057000
	         : (byte_in == 8'h6f)? 32'h6dac7000
	         : (byte_in == 8'h70)? 32'h16444000
	         : (byte_in == 8'h71)? 32'hdded4000
	         : (byte_in == 8'h72)? 32'ha9785000
	         : (byte_in == 8'h73)? 32'h62d15000
	         : (byte_in == 8'h74)? 32'h81174000
	         : (byte_in == 8'h75)? 32'h4abe4000
	         : (byte_in == 8'h76)? 32'h3e2b5000
	         : (byte_in == 8'h77)? 32'hf5825000
	         : (byte_in == 8'h78)? 32'h683d6000
	         : (byte_in == 8'h79)? 32'ha3946000
	         : (byte_in == 8'h7a)? 32'hd7017000
	         : (byte_in == 8'h7b)? 32'h1ca87000
	         : (byte_in == 8'h7c)? 32'hff6e6000
	         : (byte_in == 8'h7d)? 32'h34c76000
	         : (byte_in == 8'h7e)? 32'h40527000
	         : (byte_in == 8'h7f)? 32'h8bfb7000
	         : (byte_in == 8'h80)? 32'he0278000
	         : (byte_in == 8'h81)? 32'h2b8e8000
	         : (byte_in == 8'h82)? 32'h5f1b9000
	         : (byte_in == 8'h83)? 32'h94b29000
	         : (byte_in == 8'h84)? 32'h77748000
	         : (byte_in == 8'h85)? 32'hbcdd8000
	         : (byte_in == 8'h86)? 32'hc8489000
	         : (byte_in == 8'h87)? 32'h03e19000
	         : (byte_in == 8'h88)? 32'h9e5ea000
	         : (byte_in == 8'h89)? 32'h55f7a000
	         : (byte_in == 8'h8a)? 32'h2162b000
	         : (byte_in == 8'h8b)? 32'heacbb000
	         : (byte_in == 8'h8c)? 32'h090da000
	         : (byte_in == 8'h8d)? 32'hc2a4a000
	         : (byte_in == 8'h8e)? 32'hb631b000
	         : (byte_in == 8'h8f)? 32'h7d98b000
	         : (byte_in == 8'h90)? 32'h06708000
	         : (byte_in == 8'h91)? 32'hcdd98000
	         : (byte_in == 8'h92)? 32'hb94c9000
	         : (byte_in == 8'h93)? 32'h72e59000
	         : (byte_in == 8'h94)? 32'h91238000
	         : (byte_in == 8'h95)? 32'h5a8a8000
	         : (byte_in == 8'h96)? 32'h2e1f9000
	         : (byte_in == 8'h97)? 32'he5b69000
	         : (byte_in == 8'h98)? 32'h7809a000
	         : (byte_in == 8'h99)? 32'hb3a0a000
	         : (byte_in == 8'h9a)? 32'hc735b000
	         : (byte_in == 8'h9b)? 32'h0c9cb000
	         : (byte_in == 8'h9c)? 32'hef5aa000
	         : (byte_in == 8'h9d)? 32'h24f3a000
	         : (byte_in == 8'h9e)? 32'h5066b000
	         : (byte_in == 8'h9f)? 32'h9bcfb000
	         : (byte_in == 8'ha0)? 32'h146bc000
	         : (byte_in == 8'ha1)? 32'hdfc2c000
	         : (byte_in == 8'ha2)? 32'hab57d000
	         : (byte_in == 8'ha3)? 32'h60fed000
	         : (byte_in == 8'ha4)? 32'h8338c000
	         : (byte_in == 8'ha5)? 32'h4891c000
	         : (byte_in == 8'ha6)? 32'h3c04d000
	         : (byte_in == 8'ha7)? 32'hf7add000
	         : (byte_in == 8'ha8)? 32'h6a12e000
	         : (byte_in == 8'ha9)? 32'ha1bbe000
	         : (byte_in == 8'haa)? 32'hd52ef000
	         : (byte_in == 8'hab)? 32'h1e87f000
	         : (byte_in == 8'hac)? 32'hfd41e000
	         : (byte_in == 8'had)? 32'h36e8e000
	         : (byte_in == 8'hae)? 32'h427df000
	         : (byte_in == 8'haf)? 32'h89d4f000
	         : (byte_in == 8'hb0)? 32'hf23cc000
	         : (byte_in == 8'hb1)? 32'h3995c000
	         : (byte_in == 8'hb2)? 32'h4d00d000
	         : (byte_in == 8'hb3)? 32'h86a9d000
	         : (byte_in == 8'hb4)? 32'h656fc000
	         : (byte_in == 8'hb5)? 32'haec6c000
	         : (byte_in == 8'hb6)? 32'hda53d000
	         : (byte_in == 8'hb7)? 32'h11fad000
	         : (byte_in == 8'hb8)? 32'h8c45e000
	         : (byte_in == 8'hb9)? 32'h47ece000
	         : (byte_in == 8'hba)? 32'h3379f000
	         : (byte_in == 8'hbb)? 32'hf8d0f000
	         : (byte_in == 8'hbc)? 32'h1b16e000
	         : (byte_in == 8'hbd)? 32'hd0bfe000
	         : (byte_in == 8'hbe)? 32'ha42af000
	         : (byte_in == 8'hbf)? 32'h6f83f000
	         : (byte_in == 8'hc0)? 32'he4788000
	         : (byte_in == 8'hc1)? 32'h2fd18000
	         : (byte_in == 8'hc2)? 32'h5b449000
	         : (byte_in == 8'hc3)? 32'h90ed9000
	         : (byte_in == 8'hc4)? 32'h732b8000
	         : (byte_in == 8'hc5)? 32'hb8828000
	         : (byte_in == 8'hc6)? 32'hcc179000
	         : (byte_in == 8'hc7)? 32'h07be9000
	         : (byte_in == 8'hc8)? 32'h9a01a000
	         : (byte_in == 8'hc9)? 32'h51a8a000
	         : (byte_in == 8'hca)? 32'h253db000
	         : (byte_in == 8'hcb)? 32'hee94b000
	         : (byte_in == 8'hcc)? 32'h0d52a000
	         : (byte_in == 8'hcd)? 32'hc6fba000
	         : (byte_in == 8'hce)? 32'hb26eb000
	         : (byte_in == 8'hcf)? 32'h79c7b000
	         : (byte_in == 8'hd0)? 32'h022f8000
	         : (byte_in == 8'hd1)? 32'hc9868000
	         : (byte_in == 8'hd2)? 32'hbd139000
	         : (byte_in == 8'hd3)? 32'h76ba9000
	         : (byte_in == 8'hd4)? 32'h957c8000
	         : (byte_in == 8'hd5)? 32'h5ed58000
	         : (byte_in == 8'hd6)? 32'h2a409000
	         : (byte_in == 8'hd7)? 32'he1e99000
	         : (byte_in == 8'hd8)? 32'h7c56a000
	         : (byte_in == 8'hd9)? 32'hb7ffa000
	         : (byte_in == 8'hda)? 32'hc36ab000
	         : (byte_in == 8'hdb)? 32'h08c3b000
	         : (byte_in == 8'hdc)? 32'heb05a000
	         : (byte_in == 8'hdd)? 32'h20aca000
	         : (byte_in == 8'hde)? 32'h5439b000
	         : (byte_in == 8'hdf)? 32'h9f90b000
	         : (byte_in == 8'he0)? 32'h1034c000
	         : (byte_in == 8'he1)? 32'hdb9dc000
	         : (byte_in == 8'he2)? 32'haf08d000
	         : (byte_in == 8'he3)? 32'h64a1d000
	         : (byte_in == 8'he4)? 32'h8767c000
	         : (byte_in == 8'he5)? 32'h4ccec000
	         : (byte_in == 8'he6)? 32'h385bd000
	         : (byte_in == 8'he7)? 32'hf3f2d000
	         : (byte_in == 8'he8)? 32'h6e4de000
	         : (byte_in == 8'he9)? 32'ha5e4e000
	         : (byte_in == 8'hea)? 32'hd171f000
	         : (byte_in == 8'heb)? 32'h1ad8f000
	         : (byte_in == 8'hec)? 32'hf91ee000
	         : (byte_in == 8'hed)? 32'h32b7e000
	         : (byte_in == 8'hee)? 32'h4622f000
	         : (byte_in == 8'hef)? 32'h8d8bf000
	         : (byte_in == 8'hf0)? 32'hf663c000
	         : (byte_in == 8'hf1)? 32'h3dcac000
	         : (byte_in == 8'hf2)? 32'h495fd000
	         : (byte_in == 8'hf3)? 32'h82f6d000
	         : (byte_in == 8'hf4)? 32'h6130c000
	         : (byte_in == 8'hf5)? 32'haa99c000
	         : (byte_in == 8'hf6)? 32'hde0cd000
	         : (byte_in == 8'hf7)? 32'h15a5d000
	         : (byte_in == 8'hf8)? 32'h881ae000
	         : (byte_in == 8'hf9)? 32'h43b3e000
	         : (byte_in == 8'hfa)? 32'h3726f000
	         : (byte_in == 8'hfb)? 32'hfc8ff000
	         : (byte_in == 8'hfc)? 32'h1f49e000
	         : (byte_in == 8'hfd)? 32'hd4e0e000
	         : (byte_in == 8'hfe)? 32'ha075f000
	         :                     32'h6bdcf000;

endmodule
//}}}

module TABLE20(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h0b2de782
	         : (byte_in == 8'h02)? 32'h38942792
	         : (byte_in == 8'h03)? 32'h33b9c010
	         : (byte_in == 8'h04)? 32'h25e30f14
	         : (byte_in == 8'h05)? 32'h2ecee896
	         : (byte_in == 8'h06)? 32'h1d772886
	         : (byte_in == 8'h07)? 32'h165acf04
	         : (byte_in == 8'h08)? 32'h7a04a8a7
	         : (byte_in == 8'h09)? 32'h71294f25
	         : (byte_in == 8'h0a)? 32'h42908f35
	         : (byte_in == 8'h0b)? 32'h49bd68b7
	         : (byte_in == 8'h0c)? 32'h5fe7a7b3
	         : (byte_in == 8'h0d)? 32'h54ca4031
	         : (byte_in == 8'h0e)? 32'h67738021
	         : (byte_in == 8'h0f)? 32'h6c5e67a3
	         : (byte_in == 8'h10)? 32'h40ebf9aa
	         : (byte_in == 8'h11)? 32'h4bc61e28
	         : (byte_in == 8'h12)? 32'h787fde38
	         : (byte_in == 8'h13)? 32'h735239ba
	         : (byte_in == 8'h14)? 32'h6508f6be
	         : (byte_in == 8'h15)? 32'h6e25113c
	         : (byte_in == 8'h16)? 32'h5d9cd12c
	         : (byte_in == 8'h17)? 32'h56b136ae
	         : (byte_in == 8'h18)? 32'h3aef510d
	         : (byte_in == 8'h19)? 32'h31c2b68f
	         : (byte_in == 8'h1a)? 32'h027b769f
	         : (byte_in == 8'h1b)? 32'h0956911d
	         : (byte_in == 8'h1c)? 32'h1f0c5e19
	         : (byte_in == 8'h1d)? 32'h1421b99b
	         : (byte_in == 8'h1e)? 32'h2798798b
	         : (byte_in == 8'h1f)? 32'h2cb59e09
	         : (byte_in == 8'h20)? 32'hcc9d76dd
	         : (byte_in == 8'h21)? 32'hc7b0915f
	         : (byte_in == 8'h22)? 32'hf409514f
	         : (byte_in == 8'h23)? 32'hff24b6cd
	         : (byte_in == 8'h24)? 32'he97e79c9
	         : (byte_in == 8'h25)? 32'he2539e4b
	         : (byte_in == 8'h26)? 32'hd1ea5e5b
	         : (byte_in == 8'h27)? 32'hdac7b9d9
	         : (byte_in == 8'h28)? 32'hb699de7a
	         : (byte_in == 8'h29)? 32'hbdb439f8
	         : (byte_in == 8'h2a)? 32'h8e0df9e8
	         : (byte_in == 8'h2b)? 32'h85201e6a
	         : (byte_in == 8'h2c)? 32'h937ad16e
	         : (byte_in == 8'h2d)? 32'h985736ec
	         : (byte_in == 8'h2e)? 32'habeef6fc
	         : (byte_in == 8'h2f)? 32'ha0c3117e
	         : (byte_in == 8'h30)? 32'h8c768f77
	         : (byte_in == 8'h31)? 32'h875b68f5
	         : (byte_in == 8'h32)? 32'hb4e2a8e5
	         : (byte_in == 8'h33)? 32'hbfcf4f67
	         : (byte_in == 8'h34)? 32'ha9958063
	         : (byte_in == 8'h35)? 32'ha2b867e1
	         : (byte_in == 8'h36)? 32'h9101a7f1
	         : (byte_in == 8'h37)? 32'h9a2c4073
	         : (byte_in == 8'h38)? 32'hf67227d0
	         : (byte_in == 8'h39)? 32'hfd5fc052
	         : (byte_in == 8'h3a)? 32'hcee60042
	         : (byte_in == 8'h3b)? 32'hc5cbe7c0
	         : (byte_in == 8'h3c)? 32'hd39128c4
	         : (byte_in == 8'h3d)? 32'hd8bccf46
	         : (byte_in == 8'h3e)? 32'heb050f56
	         : (byte_in == 8'h3f)? 32'he028e8d4
	         : (byte_in == 8'h40)? 32'hb26e3344
	         : (byte_in == 8'h41)? 32'hb943d4c6
	         : (byte_in == 8'h42)? 32'h8afa14d6
	         : (byte_in == 8'h43)? 32'h81d7f354
	         : (byte_in == 8'h44)? 32'h978d3c50
	         : (byte_in == 8'h45)? 32'h9ca0dbd2
	         : (byte_in == 8'h46)? 32'haf191bc2
	         : (byte_in == 8'h47)? 32'ha434fc40
	         : (byte_in == 8'h48)? 32'hc86a9be3
	         : (byte_in == 8'h49)? 32'hc3477c61
	         : (byte_in == 8'h4a)? 32'hf0febc71
	         : (byte_in == 8'h4b)? 32'hfbd35bf3
	         : (byte_in == 8'h4c)? 32'hed8994f7
	         : (byte_in == 8'h4d)? 32'he6a47375
	         : (byte_in == 8'h4e)? 32'hd51db365
	         : (byte_in == 8'h4f)? 32'hde3054e7
	         : (byte_in == 8'h50)? 32'hf285caee
	         : (byte_in == 8'h51)? 32'hf9a82d6c
	         : (byte_in == 8'h52)? 32'hca11ed7c
	         : (byte_in == 8'h53)? 32'hc13c0afe
	         : (byte_in == 8'h54)? 32'hd766c5fa
	         : (byte_in == 8'h55)? 32'hdc4b2278
	         : (byte_in == 8'h56)? 32'heff2e268
	         : (byte_in == 8'h57)? 32'he4df05ea
	         : (byte_in == 8'h58)? 32'h88816249
	         : (byte_in == 8'h59)? 32'h83ac85cb
	         : (byte_in == 8'h5a)? 32'hb01545db
	         : (byte_in == 8'h5b)? 32'hbb38a259
	         : (byte_in == 8'h5c)? 32'had626d5d
	         : (byte_in == 8'h5d)? 32'ha64f8adf
	         : (byte_in == 8'h5e)? 32'h95f64acf
	         : (byte_in == 8'h5f)? 32'h9edbad4d
	         : (byte_in == 8'h60)? 32'h7ef34599
	         : (byte_in == 8'h61)? 32'h75dea21b
	         : (byte_in == 8'h62)? 32'h4667620b
	         : (byte_in == 8'h63)? 32'h4d4a8589
	         : (byte_in == 8'h64)? 32'h5b104a8d
	         : (byte_in == 8'h65)? 32'h503dad0f
	         : (byte_in == 8'h66)? 32'h63846d1f
	         : (byte_in == 8'h67)? 32'h68a98a9d
	         : (byte_in == 8'h68)? 32'h04f7ed3e
	         : (byte_in == 8'h69)? 32'h0fda0abc
	         : (byte_in == 8'h6a)? 32'h3c63caac
	         : (byte_in == 8'h6b)? 32'h374e2d2e
	         : (byte_in == 8'h6c)? 32'h2114e22a
	         : (byte_in == 8'h6d)? 32'h2a3905a8
	         : (byte_in == 8'h6e)? 32'h1980c5b8
	         : (byte_in == 8'h6f)? 32'h12ad223a
	         : (byte_in == 8'h70)? 32'h3e18bc33
	         : (byte_in == 8'h71)? 32'h35355bb1
	         : (byte_in == 8'h72)? 32'h068c9ba1
	         : (byte_in == 8'h73)? 32'h0da17c23
	         : (byte_in == 8'h74)? 32'h1bfbb327
	         : (byte_in == 8'h75)? 32'h10d654a5
	         : (byte_in == 8'h76)? 32'h236f94b5
	         : (byte_in == 8'h77)? 32'h28427337
	         : (byte_in == 8'h78)? 32'h441c1494
	         : (byte_in == 8'h79)? 32'h4f31f316
	         : (byte_in == 8'h7a)? 32'h7c883306
	         : (byte_in == 8'h7b)? 32'h77a5d484
	         : (byte_in == 8'h7c)? 32'h61ff1b80
	         : (byte_in == 8'h7d)? 32'h6ad2fc02
	         : (byte_in == 8'h7e)? 32'h596b3c12
	         : (byte_in == 8'h7f)? 32'h5246db90
	         : (byte_in == 8'h80)? 32'h92170a39
	         : (byte_in == 8'h81)? 32'h993aedbb
	         : (byte_in == 8'h82)? 32'haa832dab
	         : (byte_in == 8'h83)? 32'ha1aeca29
	         : (byte_in == 8'h84)? 32'hb7f4052d
	         : (byte_in == 8'h85)? 32'hbcd9e2af
	         : (byte_in == 8'h86)? 32'h8f6022bf
	         : (byte_in == 8'h87)? 32'h844dc53d
	         : (byte_in == 8'h88)? 32'he813a29e
	         : (byte_in == 8'h89)? 32'he33e451c
	         : (byte_in == 8'h8a)? 32'hd087850c
	         : (byte_in == 8'h8b)? 32'hdbaa628e
	         : (byte_in == 8'h8c)? 32'hcdf0ad8a
	         : (byte_in == 8'h8d)? 32'hc6dd4a08
	         : (byte_in == 8'h8e)? 32'hf5648a18
	         : (byte_in == 8'h8f)? 32'hfe496d9a
	         : (byte_in == 8'h90)? 32'hd2fcf393
	         : (byte_in == 8'h91)? 32'hd9d11411
	         : (byte_in == 8'h92)? 32'hea68d401
	         : (byte_in == 8'h93)? 32'he1453383
	         : (byte_in == 8'h94)? 32'hf71ffc87
	         : (byte_in == 8'h95)? 32'hfc321b05
	         : (byte_in == 8'h96)? 32'hcf8bdb15
	         : (byte_in == 8'h97)? 32'hc4a63c97
	         : (byte_in == 8'h98)? 32'ha8f85b34
	         : (byte_in == 8'h99)? 32'ha3d5bcb6
	         : (byte_in == 8'h9a)? 32'h906c7ca6
	         : (byte_in == 8'h9b)? 32'h9b419b24
	         : (byte_in == 8'h9c)? 32'h8d1b5420
	         : (byte_in == 8'h9d)? 32'h8636b3a2
	         : (byte_in == 8'h9e)? 32'hb58f73b2
	         : (byte_in == 8'h9f)? 32'hbea29430
	         : (byte_in == 8'ha0)? 32'h5e8a7ce4
	         : (byte_in == 8'ha1)? 32'h55a79b66
	         : (byte_in == 8'ha2)? 32'h661e5b76
	         : (byte_in == 8'ha3)? 32'h6d33bcf4
	         : (byte_in == 8'ha4)? 32'h7b6973f0
	         : (byte_in == 8'ha5)? 32'h70449472
	         : (byte_in == 8'ha6)? 32'h43fd5462
	         : (byte_in == 8'ha7)? 32'h48d0b3e0
	         : (byte_in == 8'ha8)? 32'h248ed443
	         : (byte_in == 8'ha9)? 32'h2fa333c1
	         : (byte_in == 8'haa)? 32'h1c1af3d1
	         : (byte_in == 8'hab)? 32'h17371453
	         : (byte_in == 8'hac)? 32'h016ddb57
	         : (byte_in == 8'had)? 32'h0a403cd5
	         : (byte_in == 8'hae)? 32'h39f9fcc5
	         : (byte_in == 8'haf)? 32'h32d41b47
	         : (byte_in == 8'hb0)? 32'h1e61854e
	         : (byte_in == 8'hb1)? 32'h154c62cc
	         : (byte_in == 8'hb2)? 32'h26f5a2dc
	         : (byte_in == 8'hb3)? 32'h2dd8455e
	         : (byte_in == 8'hb4)? 32'h3b828a5a
	         : (byte_in == 8'hb5)? 32'h30af6dd8
	         : (byte_in == 8'hb6)? 32'h0316adc8
	         : (byte_in == 8'hb7)? 32'h083b4a4a
	         : (byte_in == 8'hb8)? 32'h64652de9
	         : (byte_in == 8'hb9)? 32'h6f48ca6b
	         : (byte_in == 8'hba)? 32'h5cf10a7b
	         : (byte_in == 8'hbb)? 32'h57dcedf9
	         : (byte_in == 8'hbc)? 32'h418622fd
	         : (byte_in == 8'hbd)? 32'h4aabc57f
	         : (byte_in == 8'hbe)? 32'h7912056f
	         : (byte_in == 8'hbf)? 32'h723fe2ed
	         : (byte_in == 8'hc0)? 32'h2079397d
	         : (byte_in == 8'hc1)? 32'h2b54deff
	         : (byte_in == 8'hc2)? 32'h18ed1eef
	         : (byte_in == 8'hc3)? 32'h13c0f96d
	         : (byte_in == 8'hc4)? 32'h059a3669
	         : (byte_in == 8'hc5)? 32'h0eb7d1eb
	         : (byte_in == 8'hc6)? 32'h3d0e11fb
	         : (byte_in == 8'hc7)? 32'h3623f679
	         : (byte_in == 8'hc8)? 32'h5a7d91da
	         : (byte_in == 8'hc9)? 32'h51507658
	         : (byte_in == 8'hca)? 32'h62e9b648
	         : (byte_in == 8'hcb)? 32'h69c451ca
	         : (byte_in == 8'hcc)? 32'h7f9e9ece
	         : (byte_in == 8'hcd)? 32'h74b3794c
	         : (byte_in == 8'hce)? 32'h470ab95c
	         : (byte_in == 8'hcf)? 32'h4c275ede
	         : (byte_in == 8'hd0)? 32'h6092c0d7
	         : (byte_in == 8'hd1)? 32'h6bbf2755
	         : (byte_in == 8'hd2)? 32'h5806e745
	         : (byte_in == 8'hd3)? 32'h532b00c7
	         : (byte_in == 8'hd4)? 32'h4571cfc3
	         : (byte_in == 8'hd5)? 32'h4e5c2841
	         : (byte_in == 8'hd6)? 32'h7de5e851
	         : (byte_in == 8'hd7)? 32'h76c80fd3
	         : (byte_in == 8'hd8)? 32'h1a966870
	         : (byte_in == 8'hd9)? 32'h11bb8ff2
	         : (byte_in == 8'hda)? 32'h22024fe2
	         : (byte_in == 8'hdb)? 32'h292fa860
	         : (byte_in == 8'hdc)? 32'h3f756764
	         : (byte_in == 8'hdd)? 32'h345880e6
	         : (byte_in == 8'hde)? 32'h07e140f6
	         : (byte_in == 8'hdf)? 32'h0ccca774
	         : (byte_in == 8'he0)? 32'hece44fa0
	         : (byte_in == 8'he1)? 32'he7c9a822
	         : (byte_in == 8'he2)? 32'hd4706832
	         : (byte_in == 8'he3)? 32'hdf5d8fb0
	         : (byte_in == 8'he4)? 32'hc90740b4
	         : (byte_in == 8'he5)? 32'hc22aa736
	         : (byte_in == 8'he6)? 32'hf1936726
	         : (byte_in == 8'he7)? 32'hfabe80a4
	         : (byte_in == 8'he8)? 32'h96e0e707
	         : (byte_in == 8'he9)? 32'h9dcd0085
	         : (byte_in == 8'hea)? 32'hae74c095
	         : (byte_in == 8'heb)? 32'ha5592717
	         : (byte_in == 8'hec)? 32'hb303e813
	         : (byte_in == 8'hed)? 32'hb82e0f91
	         : (byte_in == 8'hee)? 32'h8b97cf81
	         : (byte_in == 8'hef)? 32'h80ba2803
	         : (byte_in == 8'hf0)? 32'hac0fb60a
	         : (byte_in == 8'hf1)? 32'ha7225188
	         : (byte_in == 8'hf2)? 32'h949b9198
	         : (byte_in == 8'hf3)? 32'h9fb6761a
	         : (byte_in == 8'hf4)? 32'h89ecb91e
	         : (byte_in == 8'hf5)? 32'h82c15e9c
	         : (byte_in == 8'hf6)? 32'hb1789e8c
	         : (byte_in == 8'hf7)? 32'hba55790e
	         : (byte_in == 8'hf8)? 32'hd60b1ead
	         : (byte_in == 8'hf9)? 32'hdd26f92f
	         : (byte_in == 8'hfa)? 32'hee9f393f
	         : (byte_in == 8'hfb)? 32'he5b2debd
	         : (byte_in == 8'hfc)? 32'hf3e811b9
	         : (byte_in == 8'hfd)? 32'hf8c5f63b
	         : (byte_in == 8'hfe)? 32'hcb7c362b
	         :                     32'hc051d1a9;

endmodule
//}}}

module TABLE21(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h64dd6689
	         : (byte_in == 8'h02)? 32'h242e1472
	         : (byte_in == 8'h03)? 32'h40f372fb
	         : (byte_in == 8'h04)? 32'hc9bacd12
	         : (byte_in == 8'h05)? 32'had67ab9b
	         : (byte_in == 8'h06)? 32'hed94d960
	         : (byte_in == 8'h07)? 32'h8949bfe9
	         : (byte_in == 8'h08)? 32'h485d28e4
	         : (byte_in == 8'h09)? 32'h2c804e6d
	         : (byte_in == 8'h0a)? 32'h6c733c96
	         : (byte_in == 8'h0b)? 32'h08ae5a1f
	         : (byte_in == 8'h0c)? 32'h81e7e5f6
	         : (byte_in == 8'h0d)? 32'he53a837f
	         : (byte_in == 8'h0e)? 32'ha5c9f184
	         : (byte_in == 8'h0f)? 32'hc114970d
	         : (byte_in == 8'h10)? 32'ha0cd5a34
	         : (byte_in == 8'h11)? 32'hc4103cbd
	         : (byte_in == 8'h12)? 32'h84e34e46
	         : (byte_in == 8'h13)? 32'he03e28cf
	         : (byte_in == 8'h14)? 32'h69779726
	         : (byte_in == 8'h15)? 32'h0daaf1af
	         : (byte_in == 8'h16)? 32'h4d598354
	         : (byte_in == 8'h17)? 32'h2984e5dd
	         : (byte_in == 8'h18)? 32'he89072d0
	         : (byte_in == 8'h19)? 32'h8c4d1459
	         : (byte_in == 8'h1a)? 32'hccbe66a2
	         : (byte_in == 8'h1b)? 32'ha863002b
	         : (byte_in == 8'h1c)? 32'h212abfc2
	         : (byte_in == 8'h1d)? 32'h45f7d94b
	         : (byte_in == 8'h1e)? 32'h0504abb0
	         : (byte_in == 8'h1f)? 32'h61d9cd39
	         : (byte_in == 8'h20)? 32'h9b96b64a
	         : (byte_in == 8'h21)? 32'hff4bd0c3
	         : (byte_in == 8'h22)? 32'hbfb8a238
	         : (byte_in == 8'h23)? 32'hdb65c4b1
	         : (byte_in == 8'h24)? 32'h522c7b58
	         : (byte_in == 8'h25)? 32'h36f11dd1
	         : (byte_in == 8'h26)? 32'h76026f2a
	         : (byte_in == 8'h27)? 32'h12df09a3
	         : (byte_in == 8'h28)? 32'hd3cb9eae
	         : (byte_in == 8'h29)? 32'hb716f827
	         : (byte_in == 8'h2a)? 32'hf7e58adc
	         : (byte_in == 8'h2b)? 32'h9338ec55
	         : (byte_in == 8'h2c)? 32'h1a7153bc
	         : (byte_in == 8'h2d)? 32'h7eac3535
	         : (byte_in == 8'h2e)? 32'h3e5f47ce
	         : (byte_in == 8'h2f)? 32'h5a822147
	         : (byte_in == 8'h30)? 32'h3b5bec7e
	         : (byte_in == 8'h31)? 32'h5f868af7
	         : (byte_in == 8'h32)? 32'h1f75f80c
	         : (byte_in == 8'h33)? 32'h7ba89e85
	         : (byte_in == 8'h34)? 32'hf2e1216c
	         : (byte_in == 8'h35)? 32'h963c47e5
	         : (byte_in == 8'h36)? 32'hd6cf351e
	         : (byte_in == 8'h37)? 32'hb2125397
	         : (byte_in == 8'h38)? 32'h7306c49a
	         : (byte_in == 8'h39)? 32'h17dba213
	         : (byte_in == 8'h3a)? 32'h5728d0e8
	         : (byte_in == 8'h3b)? 32'h33f5b661
	         : (byte_in == 8'h3c)? 32'hbabc0988
	         : (byte_in == 8'h3d)? 32'hde616f01
	         : (byte_in == 8'h3e)? 32'h9e921dfa
	         : (byte_in == 8'h3f)? 32'hfa4f7b73
	         : (byte_in == 8'h40)? 32'h4ab753eb
	         : (byte_in == 8'h41)? 32'h2e6a3562
	         : (byte_in == 8'h42)? 32'h6e994799
	         : (byte_in == 8'h43)? 32'h0a442110
	         : (byte_in == 8'h44)? 32'h830d9ef9
	         : (byte_in == 8'h45)? 32'he7d0f870
	         : (byte_in == 8'h46)? 32'ha7238a8b
	         : (byte_in == 8'h47)? 32'hc3feec02
	         : (byte_in == 8'h48)? 32'h02ea7b0f
	         : (byte_in == 8'h49)? 32'h66371d86
	         : (byte_in == 8'h4a)? 32'h26c46f7d
	         : (byte_in == 8'h4b)? 32'h421909f4
	         : (byte_in == 8'h4c)? 32'hcb50b61d
	         : (byte_in == 8'h4d)? 32'haf8dd094
	         : (byte_in == 8'h4e)? 32'hef7ea26f
	         : (byte_in == 8'h4f)? 32'h8ba3c4e6
	         : (byte_in == 8'h50)? 32'hea7a09df
	         : (byte_in == 8'h51)? 32'h8ea76f56
	         : (byte_in == 8'h52)? 32'hce541dad
	         : (byte_in == 8'h53)? 32'haa897b24
	         : (byte_in == 8'h54)? 32'h23c0c4cd
	         : (byte_in == 8'h55)? 32'h471da244
	         : (byte_in == 8'h56)? 32'h07eed0bf
	         : (byte_in == 8'h57)? 32'h6333b636
	         : (byte_in == 8'h58)? 32'ha227213b
	         : (byte_in == 8'h59)? 32'hc6fa47b2
	         : (byte_in == 8'h5a)? 32'h86093549
	         : (byte_in == 8'h5b)? 32'he2d453c0
	         : (byte_in == 8'h5c)? 32'h6b9dec29
	         : (byte_in == 8'h5d)? 32'h0f408aa0
	         : (byte_in == 8'h5e)? 32'h4fb3f85b
	         : (byte_in == 8'h5f)? 32'h2b6e9ed2
	         : (byte_in == 8'h60)? 32'hd121e5a1
	         : (byte_in == 8'h61)? 32'hb5fc8328
	         : (byte_in == 8'h62)? 32'hf50ff1d3
	         : (byte_in == 8'h63)? 32'h91d2975a
	         : (byte_in == 8'h64)? 32'h189b28b3
	         : (byte_in == 8'h65)? 32'h7c464e3a
	         : (byte_in == 8'h66)? 32'h3cb53cc1
	         : (byte_in == 8'h67)? 32'h58685a48
	         : (byte_in == 8'h68)? 32'h997ccd45
	         : (byte_in == 8'h69)? 32'hfda1abcc
	         : (byte_in == 8'h6a)? 32'hbd52d937
	         : (byte_in == 8'h6b)? 32'hd98fbfbe
	         : (byte_in == 8'h6c)? 32'h50c60057
	         : (byte_in == 8'h6d)? 32'h341b66de
	         : (byte_in == 8'h6e)? 32'h74e81425
	         : (byte_in == 8'h6f)? 32'h103572ac
	         : (byte_in == 8'h70)? 32'h71ecbf95
	         : (byte_in == 8'h71)? 32'h1531d91c
	         : (byte_in == 8'h72)? 32'h55c2abe7
	         : (byte_in == 8'h73)? 32'h311fcd6e
	         : (byte_in == 8'h74)? 32'hb8567287
	         : (byte_in == 8'h75)? 32'hdc8b140e
	         : (byte_in == 8'h76)? 32'h9c7866f5
	         : (byte_in == 8'h77)? 32'hf8a5007c
	         : (byte_in == 8'h78)? 32'h39b19771
	         : (byte_in == 8'h79)? 32'h5d6cf1f8
	         : (byte_in == 8'h7a)? 32'h1d9f8303
	         : (byte_in == 8'h7b)? 32'h7942e58a
	         : (byte_in == 8'h7c)? 32'hf00b5a63
	         : (byte_in == 8'h7d)? 32'h94d63cea
	         : (byte_in == 8'h7e)? 32'hd4254e11
	         : (byte_in == 8'h7f)? 32'hb0f82898
	         : (byte_in == 8'h80)? 32'h0fb84b07
	         : (byte_in == 8'h81)? 32'h6b652d8e
	         : (byte_in == 8'h82)? 32'h2b965f75
	         : (byte_in == 8'h83)? 32'h4f4b39fc
	         : (byte_in == 8'h84)? 32'hc6028615
	         : (byte_in == 8'h85)? 32'ha2dfe09c
	         : (byte_in == 8'h86)? 32'he22c9267
	         : (byte_in == 8'h87)? 32'h86f1f4ee
	         : (byte_in == 8'h88)? 32'h47e563e3
	         : (byte_in == 8'h89)? 32'h2338056a
	         : (byte_in == 8'h8a)? 32'h63cb7791
	         : (byte_in == 8'h8b)? 32'h07161118
	         : (byte_in == 8'h8c)? 32'h8e5faef1
	         : (byte_in == 8'h8d)? 32'hea82c878
	         : (byte_in == 8'h8e)? 32'haa71ba83
	         : (byte_in == 8'h8f)? 32'hceacdc0a
	         : (byte_in == 8'h90)? 32'haf751133
	         : (byte_in == 8'h91)? 32'hcba877ba
	         : (byte_in == 8'h92)? 32'h8b5b0541
	         : (byte_in == 8'h93)? 32'hef8663c8
	         : (byte_in == 8'h94)? 32'h66cfdc21
	         : (byte_in == 8'h95)? 32'h0212baa8
	         : (byte_in == 8'h96)? 32'h42e1c853
	         : (byte_in == 8'h97)? 32'h263caeda
	         : (byte_in == 8'h98)? 32'he72839d7
	         : (byte_in == 8'h99)? 32'h83f55f5e
	         : (byte_in == 8'h9a)? 32'hc3062da5
	         : (byte_in == 8'h9b)? 32'ha7db4b2c
	         : (byte_in == 8'h9c)? 32'h2e92f4c5
	         : (byte_in == 8'h9d)? 32'h4a4f924c
	         : (byte_in == 8'h9e)? 32'h0abce0b7
	         : (byte_in == 8'h9f)? 32'h6e61863e
	         : (byte_in == 8'ha0)? 32'h942efd4d
	         : (byte_in == 8'ha1)? 32'hf0f39bc4
	         : (byte_in == 8'ha2)? 32'hb000e93f
	         : (byte_in == 8'ha3)? 32'hd4dd8fb6
	         : (byte_in == 8'ha4)? 32'h5d94305f
	         : (byte_in == 8'ha5)? 32'h394956d6
	         : (byte_in == 8'ha6)? 32'h79ba242d
	         : (byte_in == 8'ha7)? 32'h1d6742a4
	         : (byte_in == 8'ha8)? 32'hdc73d5a9
	         : (byte_in == 8'ha9)? 32'hb8aeb320
	         : (byte_in == 8'haa)? 32'hf85dc1db
	         : (byte_in == 8'hab)? 32'h9c80a752
	         : (byte_in == 8'hac)? 32'h15c918bb
	         : (byte_in == 8'had)? 32'h71147e32
	         : (byte_in == 8'hae)? 32'h31e70cc9
	         : (byte_in == 8'haf)? 32'h553a6a40
	         : (byte_in == 8'hb0)? 32'h34e3a779
	         : (byte_in == 8'hb1)? 32'h503ec1f0
	         : (byte_in == 8'hb2)? 32'h10cdb30b
	         : (byte_in == 8'hb3)? 32'h7410d582
	         : (byte_in == 8'hb4)? 32'hfd596a6b
	         : (byte_in == 8'hb5)? 32'h99840ce2
	         : (byte_in == 8'hb6)? 32'hd9777e19
	         : (byte_in == 8'hb7)? 32'hbdaa1890
	         : (byte_in == 8'hb8)? 32'h7cbe8f9d
	         : (byte_in == 8'hb9)? 32'h1863e914
	         : (byte_in == 8'hba)? 32'h58909bef
	         : (byte_in == 8'hbb)? 32'h3c4dfd66
	         : (byte_in == 8'hbc)? 32'hb504428f
	         : (byte_in == 8'hbd)? 32'hd1d92406
	         : (byte_in == 8'hbe)? 32'h912a56fd
	         : (byte_in == 8'hbf)? 32'hf5f73074
	         : (byte_in == 8'hc0)? 32'h450f18ec
	         : (byte_in == 8'hc1)? 32'h21d27e65
	         : (byte_in == 8'hc2)? 32'h61210c9e
	         : (byte_in == 8'hc3)? 32'h05fc6a17
	         : (byte_in == 8'hc4)? 32'h8cb5d5fe
	         : (byte_in == 8'hc5)? 32'he868b377
	         : (byte_in == 8'hc6)? 32'ha89bc18c
	         : (byte_in == 8'hc7)? 32'hcc46a705
	         : (byte_in == 8'hc8)? 32'h0d523008
	         : (byte_in == 8'hc9)? 32'h698f5681
	         : (byte_in == 8'hca)? 32'h297c247a
	         : (byte_in == 8'hcb)? 32'h4da142f3
	         : (byte_in == 8'hcc)? 32'hc4e8fd1a
	         : (byte_in == 8'hcd)? 32'ha0359b93
	         : (byte_in == 8'hce)? 32'he0c6e968
	         : (byte_in == 8'hcf)? 32'h841b8fe1
	         : (byte_in == 8'hd0)? 32'he5c242d8
	         : (byte_in == 8'hd1)? 32'h811f2451
	         : (byte_in == 8'hd2)? 32'hc1ec56aa
	         : (byte_in == 8'hd3)? 32'ha5313023
	         : (byte_in == 8'hd4)? 32'h2c788fca
	         : (byte_in == 8'hd5)? 32'h48a5e943
	         : (byte_in == 8'hd6)? 32'h08569bb8
	         : (byte_in == 8'hd7)? 32'h6c8bfd31
	         : (byte_in == 8'hd8)? 32'had9f6a3c
	         : (byte_in == 8'hd9)? 32'hc9420cb5
	         : (byte_in == 8'hda)? 32'h89b17e4e
	         : (byte_in == 8'hdb)? 32'hed6c18c7
	         : (byte_in == 8'hdc)? 32'h6425a72e
	         : (byte_in == 8'hdd)? 32'h00f8c1a7
	         : (byte_in == 8'hde)? 32'h400bb35c
	         : (byte_in == 8'hdf)? 32'h24d6d5d5
	         : (byte_in == 8'he0)? 32'hde99aea6
	         : (byte_in == 8'he1)? 32'hba44c82f
	         : (byte_in == 8'he2)? 32'hfab7bad4
	         : (byte_in == 8'he3)? 32'h9e6adc5d
	         : (byte_in == 8'he4)? 32'h172363b4
	         : (byte_in == 8'he5)? 32'h73fe053d
	         : (byte_in == 8'he6)? 32'h330d77c6
	         : (byte_in == 8'he7)? 32'h57d0114f
	         : (byte_in == 8'he8)? 32'h96c48642
	         : (byte_in == 8'he9)? 32'hf219e0cb
	         : (byte_in == 8'hea)? 32'hb2ea9230
	         : (byte_in == 8'heb)? 32'hd637f4b9
	         : (byte_in == 8'hec)? 32'h5f7e4b50
	         : (byte_in == 8'hed)? 32'h3ba32dd9
	         : (byte_in == 8'hee)? 32'h7b505f22
	         : (byte_in == 8'hef)? 32'h1f8d39ab
	         : (byte_in == 8'hf0)? 32'h7e54f492
	         : (byte_in == 8'hf1)? 32'h1a89921b
	         : (byte_in == 8'hf2)? 32'h5a7ae0e0
	         : (byte_in == 8'hf3)? 32'h3ea78669
	         : (byte_in == 8'hf4)? 32'hb7ee3980
	         : (byte_in == 8'hf5)? 32'hd3335f09
	         : (byte_in == 8'hf6)? 32'h93c02df2
	         : (byte_in == 8'hf7)? 32'hf71d4b7b
	         : (byte_in == 8'hf8)? 32'h3609dc76
	         : (byte_in == 8'hf9)? 32'h52d4baff
	         : (byte_in == 8'hfa)? 32'h1227c804
	         : (byte_in == 8'hfb)? 32'h76faae8d
	         : (byte_in == 8'hfc)? 32'hffb31164
	         : (byte_in == 8'hfd)? 32'h9b6e77ed
	         : (byte_in == 8'hfe)? 32'hdb9d0516
	         :                     32'hbf40639f;

endmodule
//}}}

module TABLE22(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h956fa7d6
	         : (byte_in == 8'h02)? 32'h1f70960e
	         : (byte_in == 8'h03)? 32'h8a1f31d8
	         : (byte_in == 8'h04)? 32'h124b683e
	         : (byte_in == 8'h05)? 32'h8724cfe8
	         : (byte_in == 8'h06)? 32'h0d3bfe30
	         : (byte_in == 8'h07)? 32'h985459e6
	         : (byte_in == 8'h08)? 32'h0d59ec0d
	         : (byte_in == 8'h09)? 32'h98364bdb
	         : (byte_in == 8'h0a)? 32'h12297a03
	         : (byte_in == 8'h0b)? 32'h8746ddd5
	         : (byte_in == 8'h0c)? 32'h1f128433
	         : (byte_in == 8'h0d)? 32'h8a7d23e5
	         : (byte_in == 8'h0e)? 32'h0062123d
	         : (byte_in == 8'h0f)? 32'h950db5eb
	         : (byte_in == 8'h10)? 32'h2fba37ff
	         : (byte_in == 8'h11)? 32'hbad59029
	         : (byte_in == 8'h12)? 32'h30caa1f1
	         : (byte_in == 8'h13)? 32'ha5a50627
	         : (byte_in == 8'h14)? 32'h3df15fc1
	         : (byte_in == 8'h15)? 32'ha89ef817
	         : (byte_in == 8'h16)? 32'h2281c9cf
	         : (byte_in == 8'h17)? 32'hb7ee6e19
	         : (byte_in == 8'h18)? 32'h22e3dbf2
	         : (byte_in == 8'h19)? 32'hb78c7c24
	         : (byte_in == 8'h1a)? 32'h3d934dfc
	         : (byte_in == 8'h1b)? 32'ha8fcea2a
	         : (byte_in == 8'h1c)? 32'h30a8b3cc
	         : (byte_in == 8'h1d)? 32'ha5c7141a
	         : (byte_in == 8'h1e)? 32'h2fd825c2
	         : (byte_in == 8'h1f)? 32'hbab78214
	         : (byte_in == 8'h20)? 32'h2227ff88
	         : (byte_in == 8'h21)? 32'hb748585e
	         : (byte_in == 8'h22)? 32'h3d576986
	         : (byte_in == 8'h23)? 32'ha838ce50
	         : (byte_in == 8'h24)? 32'h306c97b6
	         : (byte_in == 8'h25)? 32'ha5033060
	         : (byte_in == 8'h26)? 32'h2f1c01b8
	         : (byte_in == 8'h27)? 32'hba73a66e
	         : (byte_in == 8'h28)? 32'h2f7e1385
	         : (byte_in == 8'h29)? 32'hba11b453
	         : (byte_in == 8'h2a)? 32'h300e858b
	         : (byte_in == 8'h2b)? 32'ha561225d
	         : (byte_in == 8'h2c)? 32'h3d357bbb
	         : (byte_in == 8'h2d)? 32'ha85adc6d
	         : (byte_in == 8'h2e)? 32'h2245edb5
	         : (byte_in == 8'h2f)? 32'hb72a4a63
	         : (byte_in == 8'h30)? 32'h0d9dc877
	         : (byte_in == 8'h31)? 32'h98f26fa1
	         : (byte_in == 8'h32)? 32'h12ed5e79
	         : (byte_in == 8'h33)? 32'h8782f9af
	         : (byte_in == 8'h34)? 32'h1fd6a049
	         : (byte_in == 8'h35)? 32'h8ab9079f
	         : (byte_in == 8'h36)? 32'h00a63647
	         : (byte_in == 8'h37)? 32'h95c99191
	         : (byte_in == 8'h38)? 32'h00c4247a
	         : (byte_in == 8'h39)? 32'h95ab83ac
	         : (byte_in == 8'h3a)? 32'h1fb4b274
	         : (byte_in == 8'h3b)? 32'h8adb15a2
	         : (byte_in == 8'h3c)? 32'h128f4c44
	         : (byte_in == 8'h3d)? 32'h87e0eb92
	         : (byte_in == 8'h3e)? 32'h0dffda4a
	         : (byte_in == 8'h3f)? 32'h98907d9c
	         : (byte_in == 8'h40)? 32'h5459887d
	         : (byte_in == 8'h41)? 32'hc1362fab
	         : (byte_in == 8'h42)? 32'h4b291e73
	         : (byte_in == 8'h43)? 32'hde46b9a5
	         : (byte_in == 8'h44)? 32'h4612e043
	         : (byte_in == 8'h45)? 32'hd37d4795
	         : (byte_in == 8'h46)? 32'h5962764d
	         : (byte_in == 8'h47)? 32'hcc0dd19b
	         : (byte_in == 8'h48)? 32'h59006470
	         : (byte_in == 8'h49)? 32'hcc6fc3a6
	         : (byte_in == 8'h4a)? 32'h4670f27e
	         : (byte_in == 8'h4b)? 32'hd31f55a8
	         : (byte_in == 8'h4c)? 32'h4b4b0c4e
	         : (byte_in == 8'h4d)? 32'hde24ab98
	         : (byte_in == 8'h4e)? 32'h543b9a40
	         : (byte_in == 8'h4f)? 32'hc1543d96
	         : (byte_in == 8'h50)? 32'h7be3bf82
	         : (byte_in == 8'h51)? 32'hee8c1854
	         : (byte_in == 8'h52)? 32'h6493298c
	         : (byte_in == 8'h53)? 32'hf1fc8e5a
	         : (byte_in == 8'h54)? 32'h69a8d7bc
	         : (byte_in == 8'h55)? 32'hfcc7706a
	         : (byte_in == 8'h56)? 32'h76d841b2
	         : (byte_in == 8'h57)? 32'he3b7e664
	         : (byte_in == 8'h58)? 32'h76ba538f
	         : (byte_in == 8'h59)? 32'he3d5f459
	         : (byte_in == 8'h5a)? 32'h69cac581
	         : (byte_in == 8'h5b)? 32'hfca56257
	         : (byte_in == 8'h5c)? 32'h64f13bb1
	         : (byte_in == 8'h5d)? 32'hf19e9c67
	         : (byte_in == 8'h5e)? 32'h7b81adbf
	         : (byte_in == 8'h5f)? 32'heeee0a69
	         : (byte_in == 8'h60)? 32'h767e77f5
	         : (byte_in == 8'h61)? 32'he311d023
	         : (byte_in == 8'h62)? 32'h690ee1fb
	         : (byte_in == 8'h63)? 32'hfc61462d
	         : (byte_in == 8'h64)? 32'h64351fcb
	         : (byte_in == 8'h65)? 32'hf15ab81d
	         : (byte_in == 8'h66)? 32'h7b4589c5
	         : (byte_in == 8'h67)? 32'hee2a2e13
	         : (byte_in == 8'h68)? 32'h7b279bf8
	         : (byte_in == 8'h69)? 32'hee483c2e
	         : (byte_in == 8'h6a)? 32'h64570df6
	         : (byte_in == 8'h6b)? 32'hf138aa20
	         : (byte_in == 8'h6c)? 32'h696cf3c6
	         : (byte_in == 8'h6d)? 32'hfc035410
	         : (byte_in == 8'h6e)? 32'h761c65c8
	         : (byte_in == 8'h6f)? 32'he373c21e
	         : (byte_in == 8'h70)? 32'h59c4400a
	         : (byte_in == 8'h71)? 32'hccabe7dc
	         : (byte_in == 8'h72)? 32'h46b4d604
	         : (byte_in == 8'h73)? 32'hd3db71d2
	         : (byte_in == 8'h74)? 32'h4b8f2834
	         : (byte_in == 8'h75)? 32'hdee08fe2
	         : (byte_in == 8'h76)? 32'h54ffbe3a
	         : (byte_in == 8'h77)? 32'hc19019ec
	         : (byte_in == 8'h78)? 32'h549dac07
	         : (byte_in == 8'h79)? 32'hc1f20bd1
	         : (byte_in == 8'h7a)? 32'h4bed3a09
	         : (byte_in == 8'h7b)? 32'hde829ddf
	         : (byte_in == 8'h7c)? 32'h46d6c439
	         : (byte_in == 8'h7d)? 32'hd3b963ef
	         : (byte_in == 8'h7e)? 32'h59a65237
	         : (byte_in == 8'h7f)? 32'hccc9f5e1
	         : (byte_in == 8'h80)? 32'h7cdad883
	         : (byte_in == 8'h81)? 32'he9b57f55
	         : (byte_in == 8'h82)? 32'h63aa4e8d
	         : (byte_in == 8'h83)? 32'hf6c5e95b
	         : (byte_in == 8'h84)? 32'h6e91b0bd
	         : (byte_in == 8'h85)? 32'hfbfe176b
	         : (byte_in == 8'h86)? 32'h71e126b3
	         : (byte_in == 8'h87)? 32'he48e8165
	         : (byte_in == 8'h88)? 32'h7183348e
	         : (byte_in == 8'h89)? 32'he4ec9358
	         : (byte_in == 8'h8a)? 32'h6ef3a280
	         : (byte_in == 8'h8b)? 32'hfb9c0556
	         : (byte_in == 8'h8c)? 32'h63c85cb0
	         : (byte_in == 8'h8d)? 32'hf6a7fb66
	         : (byte_in == 8'h8e)? 32'h7cb8cabe
	         : (byte_in == 8'h8f)? 32'he9d76d68
	         : (byte_in == 8'h90)? 32'h5360ef7c
	         : (byte_in == 8'h91)? 32'hc60f48aa
	         : (byte_in == 8'h92)? 32'h4c107972
	         : (byte_in == 8'h93)? 32'hd97fdea4
	         : (byte_in == 8'h94)? 32'h412b8742
	         : (byte_in == 8'h95)? 32'hd4442094
	         : (byte_in == 8'h96)? 32'h5e5b114c
	         : (byte_in == 8'h97)? 32'hcb34b69a
	         : (byte_in == 8'h98)? 32'h5e390371
	         : (byte_in == 8'h99)? 32'hcb56a4a7
	         : (byte_in == 8'h9a)? 32'h4149957f
	         : (byte_in == 8'h9b)? 32'hd42632a9
	         : (byte_in == 8'h9c)? 32'h4c726b4f
	         : (byte_in == 8'h9d)? 32'hd91dcc99
	         : (byte_in == 8'h9e)? 32'h5302fd41
	         : (byte_in == 8'h9f)? 32'hc66d5a97
	         : (byte_in == 8'ha0)? 32'h5efd270b
	         : (byte_in == 8'ha1)? 32'hcb9280dd
	         : (byte_in == 8'ha2)? 32'h418db105
	         : (byte_in == 8'ha3)? 32'hd4e216d3
	         : (byte_in == 8'ha4)? 32'h4cb64f35
	         : (byte_in == 8'ha5)? 32'hd9d9e8e3
	         : (byte_in == 8'ha6)? 32'h53c6d93b
	         : (byte_in == 8'ha7)? 32'hc6a97eed
	         : (byte_in == 8'ha8)? 32'h53a4cb06
	         : (byte_in == 8'ha9)? 32'hc6cb6cd0
	         : (byte_in == 8'haa)? 32'h4cd45d08
	         : (byte_in == 8'hab)? 32'hd9bbfade
	         : (byte_in == 8'hac)? 32'h41efa338
	         : (byte_in == 8'had)? 32'hd48004ee
	         : (byte_in == 8'hae)? 32'h5e9f3536
	         : (byte_in == 8'haf)? 32'hcbf092e0
	         : (byte_in == 8'hb0)? 32'h714710f4
	         : (byte_in == 8'hb1)? 32'he428b722
	         : (byte_in == 8'hb2)? 32'h6e3786fa
	         : (byte_in == 8'hb3)? 32'hfb58212c
	         : (byte_in == 8'hb4)? 32'h630c78ca
	         : (byte_in == 8'hb5)? 32'hf663df1c
	         : (byte_in == 8'hb6)? 32'h7c7ceec4
	         : (byte_in == 8'hb7)? 32'he9134912
	         : (byte_in == 8'hb8)? 32'h7c1efcf9
	         : (byte_in == 8'hb9)? 32'he9715b2f
	         : (byte_in == 8'hba)? 32'h636e6af7
	         : (byte_in == 8'hbb)? 32'hf601cd21
	         : (byte_in == 8'hbc)? 32'h6e5594c7
	         : (byte_in == 8'hbd)? 32'hfb3a3311
	         : (byte_in == 8'hbe)? 32'h712502c9
	         : (byte_in == 8'hbf)? 32'he44aa51f
	         : (byte_in == 8'hc0)? 32'h288350fe
	         : (byte_in == 8'hc1)? 32'hbdecf728
	         : (byte_in == 8'hc2)? 32'h37f3c6f0
	         : (byte_in == 8'hc3)? 32'ha29c6126
	         : (byte_in == 8'hc4)? 32'h3ac838c0
	         : (byte_in == 8'hc5)? 32'hafa79f16
	         : (byte_in == 8'hc6)? 32'h25b8aece
	         : (byte_in == 8'hc7)? 32'hb0d70918
	         : (byte_in == 8'hc8)? 32'h25dabcf3
	         : (byte_in == 8'hc9)? 32'hb0b51b25
	         : (byte_in == 8'hca)? 32'h3aaa2afd
	         : (byte_in == 8'hcb)? 32'hafc58d2b
	         : (byte_in == 8'hcc)? 32'h3791d4cd
	         : (byte_in == 8'hcd)? 32'ha2fe731b
	         : (byte_in == 8'hce)? 32'h28e142c3
	         : (byte_in == 8'hcf)? 32'hbd8ee515
	         : (byte_in == 8'hd0)? 32'h07396701
	         : (byte_in == 8'hd1)? 32'h9256c0d7
	         : (byte_in == 8'hd2)? 32'h1849f10f
	         : (byte_in == 8'hd3)? 32'h8d2656d9
	         : (byte_in == 8'hd4)? 32'h15720f3f
	         : (byte_in == 8'hd5)? 32'h801da8e9
	         : (byte_in == 8'hd6)? 32'h0a029931
	         : (byte_in == 8'hd7)? 32'h9f6d3ee7
	         : (byte_in == 8'hd8)? 32'h0a608b0c
	         : (byte_in == 8'hd9)? 32'h9f0f2cda
	         : (byte_in == 8'hda)? 32'h15101d02
	         : (byte_in == 8'hdb)? 32'h807fbad4
	         : (byte_in == 8'hdc)? 32'h182be332
	         : (byte_in == 8'hdd)? 32'h8d4444e4
	         : (byte_in == 8'hde)? 32'h075b753c
	         : (byte_in == 8'hdf)? 32'h9234d2ea
	         : (byte_in == 8'he0)? 32'h0aa4af76
	         : (byte_in == 8'he1)? 32'h9fcb08a0
	         : (byte_in == 8'he2)? 32'h15d43978
	         : (byte_in == 8'he3)? 32'h80bb9eae
	         : (byte_in == 8'he4)? 32'h18efc748
	         : (byte_in == 8'he5)? 32'h8d80609e
	         : (byte_in == 8'he6)? 32'h079f5146
	         : (byte_in == 8'he7)? 32'h92f0f690
	         : (byte_in == 8'he8)? 32'h07fd437b
	         : (byte_in == 8'he9)? 32'h9292e4ad
	         : (byte_in == 8'hea)? 32'h188dd575
	         : (byte_in == 8'heb)? 32'h8de272a3
	         : (byte_in == 8'hec)? 32'h15b62b45
	         : (byte_in == 8'hed)? 32'h80d98c93
	         : (byte_in == 8'hee)? 32'h0ac6bd4b
	         : (byte_in == 8'hef)? 32'h9fa91a9d
	         : (byte_in == 8'hf0)? 32'h251e9889
	         : (byte_in == 8'hf1)? 32'hb0713f5f
	         : (byte_in == 8'hf2)? 32'h3a6e0e87
	         : (byte_in == 8'hf3)? 32'haf01a951
	         : (byte_in == 8'hf4)? 32'h3755f0b7
	         : (byte_in == 8'hf5)? 32'ha23a5761
	         : (byte_in == 8'hf6)? 32'h282566b9
	         : (byte_in == 8'hf7)? 32'hbd4ac16f
	         : (byte_in == 8'hf8)? 32'h28477484
	         : (byte_in == 8'hf9)? 32'hbd28d352
	         : (byte_in == 8'hfa)? 32'h3737e28a
	         : (byte_in == 8'hfb)? 32'ha258455c
	         : (byte_in == 8'hfc)? 32'h3a0c1cba
	         : (byte_in == 8'hfd)? 32'haf63bb6c
	         : (byte_in == 8'hfe)? 32'h257c8ab4
	         :                     32'hb0132d62;

endmodule
//}}}

module TABLE23(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h90273769
	         : (byte_in == 8'h02)? 32'hca0c7117
	         : (byte_in == 8'h03)? 32'h5a2b467e
	         : (byte_in == 8'h04)? 32'h204f6ed3
	         : (byte_in == 8'h05)? 32'hb06859ba
	         : (byte_in == 8'h06)? 32'hea431fc4
	         : (byte_in == 8'h07)? 32'h7a6428ad
	         : (byte_in == 8'h08)? 32'h9418e22f
	         : (byte_in == 8'h09)? 32'h043fd546
	         : (byte_in == 8'h0a)? 32'h5e149338
	         : (byte_in == 8'h0b)? 32'hce33a451
	         : (byte_in == 8'h0c)? 32'hb4578cfc
	         : (byte_in == 8'h0d)? 32'h2470bb95
	         : (byte_in == 8'h0e)? 32'h7e5bfdeb
	         : (byte_in == 8'h0f)? 32'hee7cca82
	         : (byte_in == 8'h10)? 32'h4bb33a25
	         : (byte_in == 8'h11)? 32'hdb940d4c
	         : (byte_in == 8'h12)? 32'h81bf4b32
	         : (byte_in == 8'h13)? 32'h11987c5b
	         : (byte_in == 8'h14)? 32'h6bfc54f6
	         : (byte_in == 8'h15)? 32'hfbdb639f
	         : (byte_in == 8'h16)? 32'ha1f025e1
	         : (byte_in == 8'h17)? 32'h31d71288
	         : (byte_in == 8'h18)? 32'hdfabd80a
	         : (byte_in == 8'h19)? 32'h4f8cef63
	         : (byte_in == 8'h1a)? 32'h15a7a91d
	         : (byte_in == 8'h1b)? 32'h85809e74
	         : (byte_in == 8'h1c)? 32'hffe4b6d9
	         : (byte_in == 8'h1d)? 32'h6fc381b0
	         : (byte_in == 8'h1e)? 32'h35e8c7ce
	         : (byte_in == 8'h1f)? 32'ha5cff0a7
	         : (byte_in == 8'h20)? 32'h10a4e3cd
	         : (byte_in == 8'h21)? 32'h8083d4a4
	         : (byte_in == 8'h22)? 32'hdaa892da
	         : (byte_in == 8'h23)? 32'h4a8fa5b3
	         : (byte_in == 8'h24)? 32'h30eb8d1e
	         : (byte_in == 8'h25)? 32'ha0ccba77
	         : (byte_in == 8'h26)? 32'hfae7fc09
	         : (byte_in == 8'h27)? 32'h6ac0cb60
	         : (byte_in == 8'h28)? 32'h84bc01e2
	         : (byte_in == 8'h29)? 32'h149b368b
	         : (byte_in == 8'h2a)? 32'h4eb070f5
	         : (byte_in == 8'h2b)? 32'hde97479c
	         : (byte_in == 8'h2c)? 32'ha4f36f31
	         : (byte_in == 8'h2d)? 32'h34d45858
	         : (byte_in == 8'h2e)? 32'h6eff1e26
	         : (byte_in == 8'h2f)? 32'hfed8294f
	         : (byte_in == 8'h30)? 32'h5b17d9e8
	         : (byte_in == 8'h31)? 32'hcb30ee81
	         : (byte_in == 8'h32)? 32'h911ba8ff
	         : (byte_in == 8'h33)? 32'h013c9f96
	         : (byte_in == 8'h34)? 32'h7b58b73b
	         : (byte_in == 8'h35)? 32'heb7f8052
	         : (byte_in == 8'h36)? 32'hb154c62c
	         : (byte_in == 8'h37)? 32'h2173f145
	         : (byte_in == 8'h38)? 32'hcf0f3bc7
	         : (byte_in == 8'h39)? 32'h5f280cae
	         : (byte_in == 8'h3a)? 32'h05034ad0
	         : (byte_in == 8'h3b)? 32'h95247db9
	         : (byte_in == 8'h3c)? 32'hef405514
	         : (byte_in == 8'h3d)? 32'h7f67627d
	         : (byte_in == 8'h3e)? 32'h254c2403
	         : (byte_in == 8'h3f)? 32'hb56b136a
	         : (byte_in == 8'h40)? 32'h9c4a93c9
	         : (byte_in == 8'h41)? 32'h0c6da4a0
	         : (byte_in == 8'h42)? 32'h5646e2de
	         : (byte_in == 8'h43)? 32'hc661d5b7
	         : (byte_in == 8'h44)? 32'hbc05fd1a
	         : (byte_in == 8'h45)? 32'h2c22ca73
	         : (byte_in == 8'h46)? 32'h76098c0d
	         : (byte_in == 8'h47)? 32'he62ebb64
	         : (byte_in == 8'h48)? 32'h085271e6
	         : (byte_in == 8'h49)? 32'h9875468f
	         : (byte_in == 8'h4a)? 32'hc25e00f1
	         : (byte_in == 8'h4b)? 32'h52793798
	         : (byte_in == 8'h4c)? 32'h281d1f35
	         : (byte_in == 8'h4d)? 32'hb83a285c
	         : (byte_in == 8'h4e)? 32'he2116e22
	         : (byte_in == 8'h4f)? 32'h7236594b
	         : (byte_in == 8'h50)? 32'hd7f9a9ec
	         : (byte_in == 8'h51)? 32'h47de9e85
	         : (byte_in == 8'h52)? 32'h1df5d8fb
	         : (byte_in == 8'h53)? 32'h8dd2ef92
	         : (byte_in == 8'h54)? 32'hf7b6c73f
	         : (byte_in == 8'h55)? 32'h6791f056
	         : (byte_in == 8'h56)? 32'h3dbab628
	         : (byte_in == 8'h57)? 32'had9d8141
	         : (byte_in == 8'h58)? 32'h43e14bc3
	         : (byte_in == 8'h59)? 32'hd3c67caa
	         : (byte_in == 8'h5a)? 32'h89ed3ad4
	         : (byte_in == 8'h5b)? 32'h19ca0dbd
	         : (byte_in == 8'h5c)? 32'h63ae2510
	         : (byte_in == 8'h5d)? 32'hf3891279
	         : (byte_in == 8'h5e)? 32'ha9a25407
	         : (byte_in == 8'h5f)? 32'h3985636e
	         : (byte_in == 8'h60)? 32'h8cee7004
	         : (byte_in == 8'h61)? 32'h1cc9476d
	         : (byte_in == 8'h62)? 32'h46e20113
	         : (byte_in == 8'h63)? 32'hd6c5367a
	         : (byte_in == 8'h64)? 32'haca11ed7
	         : (byte_in == 8'h65)? 32'h3c8629be
	         : (byte_in == 8'h66)? 32'h66ad6fc0
	         : (byte_in == 8'h67)? 32'hf68a58a9
	         : (byte_in == 8'h68)? 32'h18f6922b
	         : (byte_in == 8'h69)? 32'h88d1a542
	         : (byte_in == 8'h6a)? 32'hd2fae33c
	         : (byte_in == 8'h6b)? 32'h42ddd455
	         : (byte_in == 8'h6c)? 32'h38b9fcf8
	         : (byte_in == 8'h6d)? 32'ha89ecb91
	         : (byte_in == 8'h6e)? 32'hf2b58def
	         : (byte_in == 8'h6f)? 32'h6292ba86
	         : (byte_in == 8'h70)? 32'hc75d4a21
	         : (byte_in == 8'h71)? 32'h577a7d48
	         : (byte_in == 8'h72)? 32'h0d513b36
	         : (byte_in == 8'h73)? 32'h9d760c5f
	         : (byte_in == 8'h74)? 32'he71224f2
	         : (byte_in == 8'h75)? 32'h7735139b
	         : (byte_in == 8'h76)? 32'h2d1e55e5
	         : (byte_in == 8'h77)? 32'hbd39628c
	         : (byte_in == 8'h78)? 32'h5345a80e
	         : (byte_in == 8'h79)? 32'hc3629f67
	         : (byte_in == 8'h7a)? 32'h9949d919
	         : (byte_in == 8'h7b)? 32'h096eee70
	         : (byte_in == 8'h7c)? 32'h730ac6dd
	         : (byte_in == 8'h7d)? 32'he32df1b4
	         : (byte_in == 8'h7e)? 32'hb906b7ca
	         : (byte_in == 8'h7f)? 32'h292180a3
	         : (byte_in == 8'h80)? 32'h19dce008
	         : (byte_in == 8'h81)? 32'h89fbd761
	         : (byte_in == 8'h82)? 32'hd3d0911f
	         : (byte_in == 8'h83)? 32'h43f7a676
	         : (byte_in == 8'h84)? 32'h39938edb
	         : (byte_in == 8'h85)? 32'ha9b4b9b2
	         : (byte_in == 8'h86)? 32'hf39fffcc
	         : (byte_in == 8'h87)? 32'h63b8c8a5
	         : (byte_in == 8'h88)? 32'h8dc40227
	         : (byte_in == 8'h89)? 32'h1de3354e
	         : (byte_in == 8'h8a)? 32'h47c87330
	         : (byte_in == 8'h8b)? 32'hd7ef4459
	         : (byte_in == 8'h8c)? 32'had8b6cf4
	         : (byte_in == 8'h8d)? 32'h3dac5b9d
	         : (byte_in == 8'h8e)? 32'h67871de3
	         : (byte_in == 8'h8f)? 32'hf7a02a8a
	         : (byte_in == 8'h90)? 32'h526fda2d
	         : (byte_in == 8'h91)? 32'hc248ed44
	         : (byte_in == 8'h92)? 32'h9863ab3a
	         : (byte_in == 8'h93)? 32'h08449c53
	         : (byte_in == 8'h94)? 32'h7220b4fe
	         : (byte_in == 8'h95)? 32'he2078397
	         : (byte_in == 8'h96)? 32'hb82cc5e9
	         : (byte_in == 8'h97)? 32'h280bf280
	         : (byte_in == 8'h98)? 32'hc6773802
	         : (byte_in == 8'h99)? 32'h56500f6b
	         : (byte_in == 8'h9a)? 32'h0c7b4915
	         : (byte_in == 8'h9b)? 32'h9c5c7e7c
	         : (byte_in == 8'h9c)? 32'he63856d1
	         : (byte_in == 8'h9d)? 32'h761f61b8
	         : (byte_in == 8'h9e)? 32'h2c3427c6
	         : (byte_in == 8'h9f)? 32'hbc1310af
	         : (byte_in == 8'ha0)? 32'h097803c5
	         : (byte_in == 8'ha1)? 32'h995f34ac
	         : (byte_in == 8'ha2)? 32'hc37472d2
	         : (byte_in == 8'ha3)? 32'h535345bb
	         : (byte_in == 8'ha4)? 32'h29376d16
	         : (byte_in == 8'ha5)? 32'hb9105a7f
	         : (byte_in == 8'ha6)? 32'he33b1c01
	         : (byte_in == 8'ha7)? 32'h731c2b68
	         : (byte_in == 8'ha8)? 32'h9d60e1ea
	         : (byte_in == 8'ha9)? 32'h0d47d683
	         : (byte_in == 8'haa)? 32'h576c90fd
	         : (byte_in == 8'hab)? 32'hc74ba794
	         : (byte_in == 8'hac)? 32'hbd2f8f39
	         : (byte_in == 8'had)? 32'h2d08b850
	         : (byte_in == 8'hae)? 32'h7723fe2e
	         : (byte_in == 8'haf)? 32'he704c947
	         : (byte_in == 8'hb0)? 32'h42cb39e0
	         : (byte_in == 8'hb1)? 32'hd2ec0e89
	         : (byte_in == 8'hb2)? 32'h88c748f7
	         : (byte_in == 8'hb3)? 32'h18e07f9e
	         : (byte_in == 8'hb4)? 32'h62845733
	         : (byte_in == 8'hb5)? 32'hf2a3605a
	         : (byte_in == 8'hb6)? 32'ha8882624
	         : (byte_in == 8'hb7)? 32'h38af114d
	         : (byte_in == 8'hb8)? 32'hd6d3dbcf
	         : (byte_in == 8'hb9)? 32'h46f4eca6
	         : (byte_in == 8'hba)? 32'h1cdfaad8
	         : (byte_in == 8'hbb)? 32'h8cf89db1
	         : (byte_in == 8'hbc)? 32'hf69cb51c
	         : (byte_in == 8'hbd)? 32'h66bb8275
	         : (byte_in == 8'hbe)? 32'h3c90c40b
	         : (byte_in == 8'hbf)? 32'hacb7f362
	         : (byte_in == 8'hc0)? 32'h859673c1
	         : (byte_in == 8'hc1)? 32'h15b144a8
	         : (byte_in == 8'hc2)? 32'h4f9a02d6
	         : (byte_in == 8'hc3)? 32'hdfbd35bf
	         : (byte_in == 8'hc4)? 32'ha5d91d12
	         : (byte_in == 8'hc5)? 32'h35fe2a7b
	         : (byte_in == 8'hc6)? 32'h6fd56c05
	         : (byte_in == 8'hc7)? 32'hfff25b6c
	         : (byte_in == 8'hc8)? 32'h118e91ee
	         : (byte_in == 8'hc9)? 32'h81a9a687
	         : (byte_in == 8'hca)? 32'hdb82e0f9
	         : (byte_in == 8'hcb)? 32'h4ba5d790
	         : (byte_in == 8'hcc)? 32'h31c1ff3d
	         : (byte_in == 8'hcd)? 32'ha1e6c854
	         : (byte_in == 8'hce)? 32'hfbcd8e2a
	         : (byte_in == 8'hcf)? 32'h6beab943
	         : (byte_in == 8'hd0)? 32'hce2549e4
	         : (byte_in == 8'hd1)? 32'h5e027e8d
	         : (byte_in == 8'hd2)? 32'h042938f3
	         : (byte_in == 8'hd3)? 32'h940e0f9a
	         : (byte_in == 8'hd4)? 32'hee6a2737
	         : (byte_in == 8'hd5)? 32'h7e4d105e
	         : (byte_in == 8'hd6)? 32'h24665620
	         : (byte_in == 8'hd7)? 32'hb4416149
	         : (byte_in == 8'hd8)? 32'h5a3dabcb
	         : (byte_in == 8'hd9)? 32'hca1a9ca2
	         : (byte_in == 8'hda)? 32'h9031dadc
	         : (byte_in == 8'hdb)? 32'h0016edb5
	         : (byte_in == 8'hdc)? 32'h7a72c518
	         : (byte_in == 8'hdd)? 32'hea55f271
	         : (byte_in == 8'hde)? 32'hb07eb40f
	         : (byte_in == 8'hdf)? 32'h20598366
	         : (byte_in == 8'he0)? 32'h9532900c
	         : (byte_in == 8'he1)? 32'h0515a765
	         : (byte_in == 8'he2)? 32'h5f3ee11b
	         : (byte_in == 8'he3)? 32'hcf19d672
	         : (byte_in == 8'he4)? 32'hb57dfedf
	         : (byte_in == 8'he5)? 32'h255ac9b6
	         : (byte_in == 8'he6)? 32'h7f718fc8
	         : (byte_in == 8'he7)? 32'hef56b8a1
	         : (byte_in == 8'he8)? 32'h012a7223
	         : (byte_in == 8'he9)? 32'h910d454a
	         : (byte_in == 8'hea)? 32'hcb260334
	         : (byte_in == 8'heb)? 32'h5b01345d
	         : (byte_in == 8'hec)? 32'h21651cf0
	         : (byte_in == 8'hed)? 32'hb1422b99
	         : (byte_in == 8'hee)? 32'heb696de7
	         : (byte_in == 8'hef)? 32'h7b4e5a8e
	         : (byte_in == 8'hf0)? 32'hde81aa29
	         : (byte_in == 8'hf1)? 32'h4ea69d40
	         : (byte_in == 8'hf2)? 32'h148ddb3e
	         : (byte_in == 8'hf3)? 32'h84aaec57
	         : (byte_in == 8'hf4)? 32'hfecec4fa
	         : (byte_in == 8'hf5)? 32'h6ee9f393
	         : (byte_in == 8'hf6)? 32'h34c2b5ed
	         : (byte_in == 8'hf7)? 32'ha4e58284
	         : (byte_in == 8'hf8)? 32'h4a994806
	         : (byte_in == 8'hf9)? 32'hdabe7f6f
	         : (byte_in == 8'hfa)? 32'h80953911
	         : (byte_in == 8'hfb)? 32'h10b20e78
	         : (byte_in == 8'hfc)? 32'h6ad626d5
	         : (byte_in == 8'hfd)? 32'hfaf111bc
	         : (byte_in == 8'hfe)? 32'ha0da57c2
	         :                     32'h30fd60ab;

endmodule
//}}}

module TABLE24(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h6bf648a4
	         : (byte_in == 8'h02)? 32'hc5f8f3a1
	         : (byte_in == 8'h03)? 32'hae0ebb05
	         : (byte_in == 8'h04)? 32'h79e22a4c
	         : (byte_in == 8'h05)? 32'h121462e8
	         : (byte_in == 8'h06)? 32'hbc1ad9ed
	         : (byte_in == 8'h07)? 32'hd7ec9149
	         : (byte_in == 8'h08)? 32'he007afe6
	         : (byte_in == 8'h09)? 32'h8bf1e742
	         : (byte_in == 8'h0a)? 32'h25ff5c47
	         : (byte_in == 8'h0b)? 32'h4e0914e3
	         : (byte_in == 8'h0c)? 32'h99e585aa
	         : (byte_in == 8'h0d)? 32'hf213cd0e
	         : (byte_in == 8'h0e)? 32'h5c1d760b
	         : (byte_in == 8'h0f)? 32'h37eb3eaf
	         : (byte_in == 8'h10)? 32'h98321c3d
	         : (byte_in == 8'h11)? 32'hf3c45499
	         : (byte_in == 8'h12)? 32'h5dcaef9c
	         : (byte_in == 8'h13)? 32'h363ca738
	         : (byte_in == 8'h14)? 32'he1d03671
	         : (byte_in == 8'h15)? 32'h8a267ed5
	         : (byte_in == 8'h16)? 32'h2428c5d0
	         : (byte_in == 8'h17)? 32'h4fde8d74
	         : (byte_in == 8'h18)? 32'h7835b3db
	         : (byte_in == 8'h19)? 32'h13c3fb7f
	         : (byte_in == 8'h1a)? 32'hbdcd407a
	         : (byte_in == 8'h1b)? 32'hd63b08de
	         : (byte_in == 8'h1c)? 32'h01d79997
	         : (byte_in == 8'h1d)? 32'h6a21d133
	         : (byte_in == 8'h1e)? 32'hc42f6a36
	         : (byte_in == 8'h1f)? 32'hafd92292
	         : (byte_in == 8'h20)? 32'h05f7ac6d
	         : (byte_in == 8'h21)? 32'h6e01e4c9
	         : (byte_in == 8'h22)? 32'hc00f5fcc
	         : (byte_in == 8'h23)? 32'habf91768
	         : (byte_in == 8'h24)? 32'h7c158621
	         : (byte_in == 8'h25)? 32'h17e3ce85
	         : (byte_in == 8'h26)? 32'hb9ed7580
	         : (byte_in == 8'h27)? 32'hd21b3d24
	         : (byte_in == 8'h28)? 32'he5f0038b
	         : (byte_in == 8'h29)? 32'h8e064b2f
	         : (byte_in == 8'h2a)? 32'h2008f02a
	         : (byte_in == 8'h2b)? 32'h4bfeb88e
	         : (byte_in == 8'h2c)? 32'h9c1229c7
	         : (byte_in == 8'h2d)? 32'hf7e46163
	         : (byte_in == 8'h2e)? 32'h59eada66
	         : (byte_in == 8'h2f)? 32'h321c92c2
	         : (byte_in == 8'h30)? 32'h9dc5b050
	         : (byte_in == 8'h31)? 32'hf633f8f4
	         : (byte_in == 8'h32)? 32'h583d43f1
	         : (byte_in == 8'h33)? 32'h33cb0b55
	         : (byte_in == 8'h34)? 32'he4279a1c
	         : (byte_in == 8'h35)? 32'h8fd1d2b8
	         : (byte_in == 8'h36)? 32'h21df69bd
	         : (byte_in == 8'h37)? 32'h4a292119
	         : (byte_in == 8'h38)? 32'h7dc21fb6
	         : (byte_in == 8'h39)? 32'h16345712
	         : (byte_in == 8'h3a)? 32'hb83aec17
	         : (byte_in == 8'h3b)? 32'hd3cca4b3
	         : (byte_in == 8'h3c)? 32'h042035fa
	         : (byte_in == 8'h3d)? 32'h6fd67d5e
	         : (byte_in == 8'h3e)? 32'hc1d8c65b
	         : (byte_in == 8'h3f)? 32'haa2e8eff
	         : (byte_in == 8'h40)? 32'h9e6a837e
	         : (byte_in == 8'h41)? 32'hf59ccbda
	         : (byte_in == 8'h42)? 32'h5b9270df
	         : (byte_in == 8'h43)? 32'h3064387b
	         : (byte_in == 8'h44)? 32'he788a932
	         : (byte_in == 8'h45)? 32'h8c7ee196
	         : (byte_in == 8'h46)? 32'h22705a93
	         : (byte_in == 8'h47)? 32'h49861237
	         : (byte_in == 8'h48)? 32'h7e6d2c98
	         : (byte_in == 8'h49)? 32'h159b643c
	         : (byte_in == 8'h4a)? 32'hbb95df39
	         : (byte_in == 8'h4b)? 32'hd063979d
	         : (byte_in == 8'h4c)? 32'h078f06d4
	         : (byte_in == 8'h4d)? 32'h6c794e70
	         : (byte_in == 8'h4e)? 32'hc277f575
	         : (byte_in == 8'h4f)? 32'ha981bdd1
	         : (byte_in == 8'h50)? 32'h06589f43
	         : (byte_in == 8'h51)? 32'h6daed7e7
	         : (byte_in == 8'h52)? 32'hc3a06ce2
	         : (byte_in == 8'h53)? 32'ha8562446
	         : (byte_in == 8'h54)? 32'h7fbab50f
	         : (byte_in == 8'h55)? 32'h144cfdab
	         : (byte_in == 8'h56)? 32'hba4246ae
	         : (byte_in == 8'h57)? 32'hd1b40e0a
	         : (byte_in == 8'h58)? 32'he65f30a5
	         : (byte_in == 8'h59)? 32'h8da97801
	         : (byte_in == 8'h5a)? 32'h23a7c304
	         : (byte_in == 8'h5b)? 32'h48518ba0
	         : (byte_in == 8'h5c)? 32'h9fbd1ae9
	         : (byte_in == 8'h5d)? 32'hf44b524d
	         : (byte_in == 8'h5e)? 32'h5a45e948
	         : (byte_in == 8'h5f)? 32'h31b3a1ec
	         : (byte_in == 8'h60)? 32'h9b9d2f13
	         : (byte_in == 8'h61)? 32'hf06b67b7
	         : (byte_in == 8'h62)? 32'h5e65dcb2
	         : (byte_in == 8'h63)? 32'h35939416
	         : (byte_in == 8'h64)? 32'he27f055f
	         : (byte_in == 8'h65)? 32'h89894dfb
	         : (byte_in == 8'h66)? 32'h2787f6fe
	         : (byte_in == 8'h67)? 32'h4c71be5a
	         : (byte_in == 8'h68)? 32'h7b9a80f5
	         : (byte_in == 8'h69)? 32'h106cc851
	         : (byte_in == 8'h6a)? 32'hbe627354
	         : (byte_in == 8'h6b)? 32'hd5943bf0
	         : (byte_in == 8'h6c)? 32'h0278aab9
	         : (byte_in == 8'h6d)? 32'h698ee21d
	         : (byte_in == 8'h6e)? 32'hc7805918
	         : (byte_in == 8'h6f)? 32'hac7611bc
	         : (byte_in == 8'h70)? 32'h03af332e
	         : (byte_in == 8'h71)? 32'h68597b8a
	         : (byte_in == 8'h72)? 32'hc657c08f
	         : (byte_in == 8'h73)? 32'hada1882b
	         : (byte_in == 8'h74)? 32'h7a4d1962
	         : (byte_in == 8'h75)? 32'h11bb51c6
	         : (byte_in == 8'h76)? 32'hbfb5eac3
	         : (byte_in == 8'h77)? 32'hd443a267
	         : (byte_in == 8'h78)? 32'he3a89cc8
	         : (byte_in == 8'h79)? 32'h885ed46c
	         : (byte_in == 8'h7a)? 32'h26506f69
	         : (byte_in == 8'h7b)? 32'h4da627cd
	         : (byte_in == 8'h7c)? 32'h9a4ab684
	         : (byte_in == 8'h7d)? 32'hf1bcfe20
	         : (byte_in == 8'h7e)? 32'h5fb24525
	         : (byte_in == 8'h7f)? 32'h34440d81
	         : (byte_in == 8'h80)? 32'h6019107f
	         : (byte_in == 8'h81)? 32'h0bef58db
	         : (byte_in == 8'h82)? 32'ha5e1e3de
	         : (byte_in == 8'h83)? 32'hce17ab7a
	         : (byte_in == 8'h84)? 32'h19fb3a33
	         : (byte_in == 8'h85)? 32'h720d7297
	         : (byte_in == 8'h86)? 32'hdc03c992
	         : (byte_in == 8'h87)? 32'hb7f58136
	         : (byte_in == 8'h88)? 32'h801ebf99
	         : (byte_in == 8'h89)? 32'hebe8f73d
	         : (byte_in == 8'h8a)? 32'h45e64c38
	         : (byte_in == 8'h8b)? 32'h2e10049c
	         : (byte_in == 8'h8c)? 32'hf9fc95d5
	         : (byte_in == 8'h8d)? 32'h920add71
	         : (byte_in == 8'h8e)? 32'h3c046674
	         : (byte_in == 8'h8f)? 32'h57f22ed0
	         : (byte_in == 8'h90)? 32'hf82b0c42
	         : (byte_in == 8'h91)? 32'h93dd44e6
	         : (byte_in == 8'h92)? 32'h3dd3ffe3
	         : (byte_in == 8'h93)? 32'h5625b747
	         : (byte_in == 8'h94)? 32'h81c9260e
	         : (byte_in == 8'h95)? 32'hea3f6eaa
	         : (byte_in == 8'h96)? 32'h4431d5af
	         : (byte_in == 8'h97)? 32'h2fc79d0b
	         : (byte_in == 8'h98)? 32'h182ca3a4
	         : (byte_in == 8'h99)? 32'h73daeb00
	         : (byte_in == 8'h9a)? 32'hddd45005
	         : (byte_in == 8'h9b)? 32'hb62218a1
	         : (byte_in == 8'h9c)? 32'h61ce89e8
	         : (byte_in == 8'h9d)? 32'h0a38c14c
	         : (byte_in == 8'h9e)? 32'ha4367a49
	         : (byte_in == 8'h9f)? 32'hcfc032ed
	         : (byte_in == 8'ha0)? 32'h65eebc12
	         : (byte_in == 8'ha1)? 32'h0e18f4b6
	         : (byte_in == 8'ha2)? 32'ha0164fb3
	         : (byte_in == 8'ha3)? 32'hcbe00717
	         : (byte_in == 8'ha4)? 32'h1c0c965e
	         : (byte_in == 8'ha5)? 32'h77fadefa
	         : (byte_in == 8'ha6)? 32'hd9f465ff
	         : (byte_in == 8'ha7)? 32'hb2022d5b
	         : (byte_in == 8'ha8)? 32'h85e913f4
	         : (byte_in == 8'ha9)? 32'hee1f5b50
	         : (byte_in == 8'haa)? 32'h4011e055
	         : (byte_in == 8'hab)? 32'h2be7a8f1
	         : (byte_in == 8'hac)? 32'hfc0b39b8
	         : (byte_in == 8'had)? 32'h97fd711c
	         : (byte_in == 8'hae)? 32'h39f3ca19
	         : (byte_in == 8'haf)? 32'h520582bd
	         : (byte_in == 8'hb0)? 32'hfddca02f
	         : (byte_in == 8'hb1)? 32'h962ae88b
	         : (byte_in == 8'hb2)? 32'h3824538e
	         : (byte_in == 8'hb3)? 32'h53d21b2a
	         : (byte_in == 8'hb4)? 32'h843e8a63
	         : (byte_in == 8'hb5)? 32'hefc8c2c7
	         : (byte_in == 8'hb6)? 32'h41c679c2
	         : (byte_in == 8'hb7)? 32'h2a303166
	         : (byte_in == 8'hb8)? 32'h1ddb0fc9
	         : (byte_in == 8'hb9)? 32'h762d476d
	         : (byte_in == 8'hba)? 32'hd823fc68
	         : (byte_in == 8'hbb)? 32'hb3d5b4cc
	         : (byte_in == 8'hbc)? 32'h64392585
	         : (byte_in == 8'hbd)? 32'h0fcf6d21
	         : (byte_in == 8'hbe)? 32'ha1c1d624
	         : (byte_in == 8'hbf)? 32'hca379e80
	         : (byte_in == 8'hc0)? 32'hfe739301
	         : (byte_in == 8'hc1)? 32'h9585dba5
	         : (byte_in == 8'hc2)? 32'h3b8b60a0
	         : (byte_in == 8'hc3)? 32'h507d2804
	         : (byte_in == 8'hc4)? 32'h8791b94d
	         : (byte_in == 8'hc5)? 32'hec67f1e9
	         : (byte_in == 8'hc6)? 32'h42694aec
	         : (byte_in == 8'hc7)? 32'h299f0248
	         : (byte_in == 8'hc8)? 32'h1e743ce7
	         : (byte_in == 8'hc9)? 32'h75827443
	         : (byte_in == 8'hca)? 32'hdb8ccf46
	         : (byte_in == 8'hcb)? 32'hb07a87e2
	         : (byte_in == 8'hcc)? 32'h679616ab
	         : (byte_in == 8'hcd)? 32'h0c605e0f
	         : (byte_in == 8'hce)? 32'ha26ee50a
	         : (byte_in == 8'hcf)? 32'hc998adae
	         : (byte_in == 8'hd0)? 32'h66418f3c
	         : (byte_in == 8'hd1)? 32'h0db7c798
	         : (byte_in == 8'hd2)? 32'ha3b97c9d
	         : (byte_in == 8'hd3)? 32'hc84f3439
	         : (byte_in == 8'hd4)? 32'h1fa3a570
	         : (byte_in == 8'hd5)? 32'h7455edd4
	         : (byte_in == 8'hd6)? 32'hda5b56d1
	         : (byte_in == 8'hd7)? 32'hb1ad1e75
	         : (byte_in == 8'hd8)? 32'h864620da
	         : (byte_in == 8'hd9)? 32'hedb0687e
	         : (byte_in == 8'hda)? 32'h43bed37b
	         : (byte_in == 8'hdb)? 32'h28489bdf
	         : (byte_in == 8'hdc)? 32'hffa40a96
	         : (byte_in == 8'hdd)? 32'h94524232
	         : (byte_in == 8'hde)? 32'h3a5cf937
	         : (byte_in == 8'hdf)? 32'h51aab193
	         : (byte_in == 8'he0)? 32'hfb843f6c
	         : (byte_in == 8'he1)? 32'h907277c8
	         : (byte_in == 8'he2)? 32'h3e7ccccd
	         : (byte_in == 8'he3)? 32'h558a8469
	         : (byte_in == 8'he4)? 32'h82661520
	         : (byte_in == 8'he5)? 32'he9905d84
	         : (byte_in == 8'he6)? 32'h479ee681
	         : (byte_in == 8'he7)? 32'h2c68ae25
	         : (byte_in == 8'he8)? 32'h1b83908a
	         : (byte_in == 8'he9)? 32'h7075d82e
	         : (byte_in == 8'hea)? 32'hde7b632b
	         : (byte_in == 8'heb)? 32'hb58d2b8f
	         : (byte_in == 8'hec)? 32'h6261bac6
	         : (byte_in == 8'hed)? 32'h0997f262
	         : (byte_in == 8'hee)? 32'ha7994967
	         : (byte_in == 8'hef)? 32'hcc6f01c3
	         : (byte_in == 8'hf0)? 32'h63b62351
	         : (byte_in == 8'hf1)? 32'h08406bf5
	         : (byte_in == 8'hf2)? 32'ha64ed0f0
	         : (byte_in == 8'hf3)? 32'hcdb89854
	         : (byte_in == 8'hf4)? 32'h1a54091d
	         : (byte_in == 8'hf5)? 32'h71a241b9
	         : (byte_in == 8'hf6)? 32'hdfacfabc
	         : (byte_in == 8'hf7)? 32'hb45ab218
	         : (byte_in == 8'hf8)? 32'h83b18cb7
	         : (byte_in == 8'hf9)? 32'he847c413
	         : (byte_in == 8'hfa)? 32'h46497f16
	         : (byte_in == 8'hfb)? 32'h2dbf37b2
	         : (byte_in == 8'hfc)? 32'hfa53a6fb
	         : (byte_in == 8'hfd)? 32'h91a5ee5f
	         : (byte_in == 8'hfe)? 32'h3fab555a
	         :                     32'h545d1dfe;

endmodule
//}}}

module TABLE25(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h3cd406fc
	         : (byte_in == 8'h02)? 32'hc03320fe
	         : (byte_in == 8'h03)? 32'hfce72602
	         : (byte_in == 8'h04)? 32'h79a90df9
	         : (byte_in == 8'h05)? 32'h457d0b05
	         : (byte_in == 8'h06)? 32'hb99a2d07
	         : (byte_in == 8'h07)? 32'h854e2bfb
	         : (byte_in == 8'h08)? 32'h806741fd
	         : (byte_in == 8'h09)? 32'hbcb34701
	         : (byte_in == 8'h0a)? 32'h40546103
	         : (byte_in == 8'h0b)? 32'h7c8067ff
	         : (byte_in == 8'h0c)? 32'hf9ce4c04
	         : (byte_in == 8'h0d)? 32'hc51a4af8
	         : (byte_in == 8'h0e)? 32'h39fd6cfa
	         : (byte_in == 8'h0f)? 32'h05296a06
	         : (byte_in == 8'h10)? 32'h5d5ca0f7
	         : (byte_in == 8'h11)? 32'h6188a60b
	         : (byte_in == 8'h12)? 32'h9d6f8009
	         : (byte_in == 8'h13)? 32'ha1bb86f5
	         : (byte_in == 8'h14)? 32'h24f5ad0e
	         : (byte_in == 8'h15)? 32'h1821abf2
	         : (byte_in == 8'h16)? 32'he4c68df0
	         : (byte_in == 8'h17)? 32'hd8128b0c
	         : (byte_in == 8'h18)? 32'hdd3be10a
	         : (byte_in == 8'h19)? 32'he1efe7f6
	         : (byte_in == 8'h1a)? 32'h1d08c1f4
	         : (byte_in == 8'h1b)? 32'h21dcc708
	         : (byte_in == 8'h1c)? 32'ha492ecf3
	         : (byte_in == 8'h1d)? 32'h9846ea0f
	         : (byte_in == 8'h1e)? 32'h64a1cc0d
	         : (byte_in == 8'h1f)? 32'h5875caf1
	         : (byte_in == 8'h20)? 32'h6b39cb5f
	         : (byte_in == 8'h21)? 32'h57edcda3
	         : (byte_in == 8'h22)? 32'hab0aeba1
	         : (byte_in == 8'h23)? 32'h97deed5d
	         : (byte_in == 8'h24)? 32'h1290c6a6
	         : (byte_in == 8'h25)? 32'h2e44c05a
	         : (byte_in == 8'h26)? 32'hd2a3e658
	         : (byte_in == 8'h27)? 32'hee77e0a4
	         : (byte_in == 8'h28)? 32'heb5e8aa2
	         : (byte_in == 8'h29)? 32'hd78a8c5e
	         : (byte_in == 8'h2a)? 32'h2b6daa5c
	         : (byte_in == 8'h2b)? 32'h17b9aca0
	         : (byte_in == 8'h2c)? 32'h92f7875b
	         : (byte_in == 8'h2d)? 32'hae2381a7
	         : (byte_in == 8'h2e)? 32'h52c4a7a5
	         : (byte_in == 8'h2f)? 32'h6e10a159
	         : (byte_in == 8'h30)? 32'h36656ba8
	         : (byte_in == 8'h31)? 32'h0ab16d54
	         : (byte_in == 8'h32)? 32'hf6564b56
	         : (byte_in == 8'h33)? 32'hca824daa
	         : (byte_in == 8'h34)? 32'h4fcc6651
	         : (byte_in == 8'h35)? 32'h731860ad
	         : (byte_in == 8'h36)? 32'h8fff46af
	         : (byte_in == 8'h37)? 32'hb32b4053
	         : (byte_in == 8'h38)? 32'hb6022a55
	         : (byte_in == 8'h39)? 32'h8ad62ca9
	         : (byte_in == 8'h3a)? 32'h76310aab
	         : (byte_in == 8'h3b)? 32'h4ae50c57
	         : (byte_in == 8'h3c)? 32'hcfab27ac
	         : (byte_in == 8'h3d)? 32'hf37f2150
	         : (byte_in == 8'h3e)? 32'h0f980752
	         : (byte_in == 8'h3f)? 32'h334c01ae
	         : (byte_in == 8'h40)? 32'hd14e094b
	         : (byte_in == 8'h41)? 32'hed9a0fb7
	         : (byte_in == 8'h42)? 32'h117d29b5
	         : (byte_in == 8'h43)? 32'h2da92f49
	         : (byte_in == 8'h44)? 32'ha8e704b2
	         : (byte_in == 8'h45)? 32'h9433024e
	         : (byte_in == 8'h46)? 32'h68d4244c
	         : (byte_in == 8'h47)? 32'h540022b0
	         : (byte_in == 8'h48)? 32'h512948b6
	         : (byte_in == 8'h49)? 32'h6dfd4e4a
	         : (byte_in == 8'h4a)? 32'h911a6848
	         : (byte_in == 8'h4b)? 32'hadce6eb4
	         : (byte_in == 8'h4c)? 32'h2880454f
	         : (byte_in == 8'h4d)? 32'h145443b3
	         : (byte_in == 8'h4e)? 32'he8b365b1
	         : (byte_in == 8'h4f)? 32'hd467634d
	         : (byte_in == 8'h50)? 32'h8c12a9bc
	         : (byte_in == 8'h51)? 32'hb0c6af40
	         : (byte_in == 8'h52)? 32'h4c218942
	         : (byte_in == 8'h53)? 32'h70f58fbe
	         : (byte_in == 8'h54)? 32'hf5bba445
	         : (byte_in == 8'h55)? 32'hc96fa2b9
	         : (byte_in == 8'h56)? 32'h358884bb
	         : (byte_in == 8'h57)? 32'h095c8247
	         : (byte_in == 8'h58)? 32'h0c75e841
	         : (byte_in == 8'h59)? 32'h30a1eebd
	         : (byte_in == 8'h5a)? 32'hcc46c8bf
	         : (byte_in == 8'h5b)? 32'hf092ce43
	         : (byte_in == 8'h5c)? 32'h75dce5b8
	         : (byte_in == 8'h5d)? 32'h4908e344
	         : (byte_in == 8'h5e)? 32'hb5efc546
	         : (byte_in == 8'h5f)? 32'h893bc3ba
	         : (byte_in == 8'h60)? 32'hba77c214
	         : (byte_in == 8'h61)? 32'h86a3c4e8
	         : (byte_in == 8'h62)? 32'h7a44e2ea
	         : (byte_in == 8'h63)? 32'h4690e416
	         : (byte_in == 8'h64)? 32'hc3decfed
	         : (byte_in == 8'h65)? 32'hff0ac911
	         : (byte_in == 8'h66)? 32'h03edef13
	         : (byte_in == 8'h67)? 32'h3f39e9ef
	         : (byte_in == 8'h68)? 32'h3a1083e9
	         : (byte_in == 8'h69)? 32'h06c48515
	         : (byte_in == 8'h6a)? 32'hfa23a317
	         : (byte_in == 8'h6b)? 32'hc6f7a5eb
	         : (byte_in == 8'h6c)? 32'h43b98e10
	         : (byte_in == 8'h6d)? 32'h7f6d88ec
	         : (byte_in == 8'h6e)? 32'h838aaeee
	         : (byte_in == 8'h6f)? 32'hbf5ea812
	         : (byte_in == 8'h70)? 32'he72b62e3
	         : (byte_in == 8'h71)? 32'hdbff641f
	         : (byte_in == 8'h72)? 32'h2718421d
	         : (byte_in == 8'h73)? 32'h1bcc44e1
	         : (byte_in == 8'h74)? 32'h9e826f1a
	         : (byte_in == 8'h75)? 32'ha25669e6
	         : (byte_in == 8'h76)? 32'h5eb14fe4
	         : (byte_in == 8'h77)? 32'h62654918
	         : (byte_in == 8'h78)? 32'h674c231e
	         : (byte_in == 8'h79)? 32'h5b9825e2
	         : (byte_in == 8'h7a)? 32'ha77f03e0
	         : (byte_in == 8'h7b)? 32'h9bab051c
	         : (byte_in == 8'h7c)? 32'h1ee52ee7
	         : (byte_in == 8'h7d)? 32'h2231281b
	         : (byte_in == 8'h7e)? 32'hded60e19
	         : (byte_in == 8'h7f)? 32'he20208e5
	         : (byte_in == 8'h80)? 32'h138a651e
	         : (byte_in == 8'h81)? 32'h2f5e63e2
	         : (byte_in == 8'h82)? 32'hd3b945e0
	         : (byte_in == 8'h83)? 32'hef6d431c
	         : (byte_in == 8'h84)? 32'h6a2368e7
	         : (byte_in == 8'h85)? 32'h56f76e1b
	         : (byte_in == 8'h86)? 32'haa104819
	         : (byte_in == 8'h87)? 32'h96c44ee5
	         : (byte_in == 8'h88)? 32'h93ed24e3
	         : (byte_in == 8'h89)? 32'haf39221f
	         : (byte_in == 8'h8a)? 32'h53de041d
	         : (byte_in == 8'h8b)? 32'h6f0a02e1
	         : (byte_in == 8'h8c)? 32'hea44291a
	         : (byte_in == 8'h8d)? 32'hd6902fe6
	         : (byte_in == 8'h8e)? 32'h2a7709e4
	         : (byte_in == 8'h8f)? 32'h16a30f18
	         : (byte_in == 8'h90)? 32'h4ed6c5e9
	         : (byte_in == 8'h91)? 32'h7202c315
	         : (byte_in == 8'h92)? 32'h8ee5e517
	         : (byte_in == 8'h93)? 32'hb231e3eb
	         : (byte_in == 8'h94)? 32'h377fc810
	         : (byte_in == 8'h95)? 32'h0babceec
	         : (byte_in == 8'h96)? 32'hf74ce8ee
	         : (byte_in == 8'h97)? 32'hcb98ee12
	         : (byte_in == 8'h98)? 32'hceb18414
	         : (byte_in == 8'h99)? 32'hf26582e8
	         : (byte_in == 8'h9a)? 32'h0e82a4ea
	         : (byte_in == 8'h9b)? 32'h3256a216
	         : (byte_in == 8'h9c)? 32'hb71889ed
	         : (byte_in == 8'h9d)? 32'h8bcc8f11
	         : (byte_in == 8'h9e)? 32'h772ba913
	         : (byte_in == 8'h9f)? 32'h4bffafef
	         : (byte_in == 8'ha0)? 32'h78b3ae41
	         : (byte_in == 8'ha1)? 32'h4467a8bd
	         : (byte_in == 8'ha2)? 32'hb8808ebf
	         : (byte_in == 8'ha3)? 32'h84548843
	         : (byte_in == 8'ha4)? 32'h011aa3b8
	         : (byte_in == 8'ha5)? 32'h3dcea544
	         : (byte_in == 8'ha6)? 32'hc1298346
	         : (byte_in == 8'ha7)? 32'hfdfd85ba
	         : (byte_in == 8'ha8)? 32'hf8d4efbc
	         : (byte_in == 8'ha9)? 32'hc400e940
	         : (byte_in == 8'haa)? 32'h38e7cf42
	         : (byte_in == 8'hab)? 32'h0433c9be
	         : (byte_in == 8'hac)? 32'h817de245
	         : (byte_in == 8'had)? 32'hbda9e4b9
	         : (byte_in == 8'hae)? 32'h414ec2bb
	         : (byte_in == 8'haf)? 32'h7d9ac447
	         : (byte_in == 8'hb0)? 32'h25ef0eb6
	         : (byte_in == 8'hb1)? 32'h193b084a
	         : (byte_in == 8'hb2)? 32'he5dc2e48
	         : (byte_in == 8'hb3)? 32'hd90828b4
	         : (byte_in == 8'hb4)? 32'h5c46034f
	         : (byte_in == 8'hb5)? 32'h609205b3
	         : (byte_in == 8'hb6)? 32'h9c7523b1
	         : (byte_in == 8'hb7)? 32'ha0a1254d
	         : (byte_in == 8'hb8)? 32'ha5884f4b
	         : (byte_in == 8'hb9)? 32'h995c49b7
	         : (byte_in == 8'hba)? 32'h65bb6fb5
	         : (byte_in == 8'hbb)? 32'h596f6949
	         : (byte_in == 8'hbc)? 32'hdc2142b2
	         : (byte_in == 8'hbd)? 32'he0f5444e
	         : (byte_in == 8'hbe)? 32'h1c12624c
	         : (byte_in == 8'hbf)? 32'h20c664b0
	         : (byte_in == 8'hc0)? 32'hc2c46c55
	         : (byte_in == 8'hc1)? 32'hfe106aa9
	         : (byte_in == 8'hc2)? 32'h02f74cab
	         : (byte_in == 8'hc3)? 32'h3e234a57
	         : (byte_in == 8'hc4)? 32'hbb6d61ac
	         : (byte_in == 8'hc5)? 32'h87b96750
	         : (byte_in == 8'hc6)? 32'h7b5e4152
	         : (byte_in == 8'hc7)? 32'h478a47ae
	         : (byte_in == 8'hc8)? 32'h42a32da8
	         : (byte_in == 8'hc9)? 32'h7e772b54
	         : (byte_in == 8'hca)? 32'h82900d56
	         : (byte_in == 8'hcb)? 32'hbe440baa
	         : (byte_in == 8'hcc)? 32'h3b0a2051
	         : (byte_in == 8'hcd)? 32'h07de26ad
	         : (byte_in == 8'hce)? 32'hfb3900af
	         : (byte_in == 8'hcf)? 32'hc7ed0653
	         : (byte_in == 8'hd0)? 32'h9f98cca2
	         : (byte_in == 8'hd1)? 32'ha34cca5e
	         : (byte_in == 8'hd2)? 32'h5fabec5c
	         : (byte_in == 8'hd3)? 32'h637feaa0
	         : (byte_in == 8'hd4)? 32'he631c15b
	         : (byte_in == 8'hd5)? 32'hdae5c7a7
	         : (byte_in == 8'hd6)? 32'h2602e1a5
	         : (byte_in == 8'hd7)? 32'h1ad6e759
	         : (byte_in == 8'hd8)? 32'h1fff8d5f
	         : (byte_in == 8'hd9)? 32'h232b8ba3
	         : (byte_in == 8'hda)? 32'hdfccada1
	         : (byte_in == 8'hdb)? 32'he318ab5d
	         : (byte_in == 8'hdc)? 32'h665680a6
	         : (byte_in == 8'hdd)? 32'h5a82865a
	         : (byte_in == 8'hde)? 32'ha665a058
	         : (byte_in == 8'hdf)? 32'h9ab1a6a4
	         : (byte_in == 8'he0)? 32'ha9fda70a
	         : (byte_in == 8'he1)? 32'h9529a1f6
	         : (byte_in == 8'he2)? 32'h69ce87f4
	         : (byte_in == 8'he3)? 32'h551a8108
	         : (byte_in == 8'he4)? 32'hd054aaf3
	         : (byte_in == 8'he5)? 32'hec80ac0f
	         : (byte_in == 8'he6)? 32'h10678a0d
	         : (byte_in == 8'he7)? 32'h2cb38cf1
	         : (byte_in == 8'he8)? 32'h299ae6f7
	         : (byte_in == 8'he9)? 32'h154ee00b
	         : (byte_in == 8'hea)? 32'he9a9c609
	         : (byte_in == 8'heb)? 32'hd57dc0f5
	         : (byte_in == 8'hec)? 32'h5033eb0e
	         : (byte_in == 8'hed)? 32'h6ce7edf2
	         : (byte_in == 8'hee)? 32'h9000cbf0
	         : (byte_in == 8'hef)? 32'hacd4cd0c
	         : (byte_in == 8'hf0)? 32'hf4a107fd
	         : (byte_in == 8'hf1)? 32'hc8750101
	         : (byte_in == 8'hf2)? 32'h34922703
	         : (byte_in == 8'hf3)? 32'h084621ff
	         : (byte_in == 8'hf4)? 32'h8d080a04
	         : (byte_in == 8'hf5)? 32'hb1dc0cf8
	         : (byte_in == 8'hf6)? 32'h4d3b2afa
	         : (byte_in == 8'hf7)? 32'h71ef2c06
	         : (byte_in == 8'hf8)? 32'h74c64600
	         : (byte_in == 8'hf9)? 32'h481240fc
	         : (byte_in == 8'hfa)? 32'hb4f566fe
	         : (byte_in == 8'hfb)? 32'h88216002
	         : (byte_in == 8'hfc)? 32'h0d6f4bf9
	         : (byte_in == 8'hfd)? 32'h31bb4d05
	         : (byte_in == 8'hfe)? 32'hcd5c6b07
	         :                     32'hf1886dfb;

endmodule
//}}}

module TABLE26(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'ha29d1297
	         : (byte_in == 8'h02)? 32'h2714ca3c
	         : (byte_in == 8'h03)? 32'h8589d8ab
	         : (byte_in == 8'h04)? 32'h80c2d68f
	         : (byte_in == 8'h05)? 32'h225fc418
	         : (byte_in == 8'h06)? 32'ha7d61cb3
	         : (byte_in == 8'h07)? 32'h054b0e24
	         : (byte_in == 8'h08)? 32'he0272f7d
	         : (byte_in == 8'h09)? 32'h42ba3dea
	         : (byte_in == 8'h0a)? 32'hc733e541
	         : (byte_in == 8'h0b)? 32'h65aef7d6
	         : (byte_in == 8'h0c)? 32'h60e5f9f2
	         : (byte_in == 8'h0d)? 32'hc278eb65
	         : (byte_in == 8'h0e)? 32'h47f133ce
	         : (byte_in == 8'h0f)? 32'he56c2159
	         : (byte_in == 8'h10)? 32'h6a72e5bb
	         : (byte_in == 8'h11)? 32'hc8eff72c
	         : (byte_in == 8'h12)? 32'h4d662f87
	         : (byte_in == 8'h13)? 32'heffb3d10
	         : (byte_in == 8'h14)? 32'heab03334
	         : (byte_in == 8'h15)? 32'h482d21a3
	         : (byte_in == 8'h16)? 32'hcda4f908
	         : (byte_in == 8'h17)? 32'h6f39eb9f
	         : (byte_in == 8'h18)? 32'h8a55cac6
	         : (byte_in == 8'h19)? 32'h28c8d851
	         : (byte_in == 8'h1a)? 32'had4100fa
	         : (byte_in == 8'h1b)? 32'h0fdc126d
	         : (byte_in == 8'h1c)? 32'h0a971c49
	         : (byte_in == 8'h1d)? 32'ha80a0ede
	         : (byte_in == 8'h1e)? 32'h2d83d675
	         : (byte_in == 8'h1f)? 32'h8f1ec4e2
	         : (byte_in == 8'h20)? 32'h05b7ad5a
	         : (byte_in == 8'h21)? 32'ha72abfcd
	         : (byte_in == 8'h22)? 32'h22a36766
	         : (byte_in == 8'h23)? 32'h803e75f1
	         : (byte_in == 8'h24)? 32'h85757bd5
	         : (byte_in == 8'h25)? 32'h27e86942
	         : (byte_in == 8'h26)? 32'ha261b1e9
	         : (byte_in == 8'h27)? 32'h00fca37e
	         : (byte_in == 8'h28)? 32'he5908227
	         : (byte_in == 8'h29)? 32'h470d90b0
	         : (byte_in == 8'h2a)? 32'hc284481b
	         : (byte_in == 8'h2b)? 32'h60195a8c
	         : (byte_in == 8'h2c)? 32'h655254a8
	         : (byte_in == 8'h2d)? 32'hc7cf463f
	         : (byte_in == 8'h2e)? 32'h42469e94
	         : (byte_in == 8'h2f)? 32'he0db8c03
	         : (byte_in == 8'h30)? 32'h6fc548e1
	         : (byte_in == 8'h31)? 32'hcd585a76
	         : (byte_in == 8'h32)? 32'h48d182dd
	         : (byte_in == 8'h33)? 32'hea4c904a
	         : (byte_in == 8'h34)? 32'hef079e6e
	         : (byte_in == 8'h35)? 32'h4d9a8cf9
	         : (byte_in == 8'h36)? 32'hc8135452
	         : (byte_in == 8'h37)? 32'h6a8e46c5
	         : (byte_in == 8'h38)? 32'h8fe2679c
	         : (byte_in == 8'h39)? 32'h2d7f750b
	         : (byte_in == 8'h3a)? 32'ha8f6ada0
	         : (byte_in == 8'h3b)? 32'h0a6bbf37
	         : (byte_in == 8'h3c)? 32'h0f20b113
	         : (byte_in == 8'h3d)? 32'hadbda384
	         : (byte_in == 8'h3e)? 32'h28347b2f
	         : (byte_in == 8'h3f)? 32'h8aa969b8
	         : (byte_in == 8'h40)? 32'hbf1283d3
	         : (byte_in == 8'h41)? 32'h1d8f9144
	         : (byte_in == 8'h42)? 32'h980649ef
	         : (byte_in == 8'h43)? 32'h3a9b5b78
	         : (byte_in == 8'h44)? 32'h3fd0555c
	         : (byte_in == 8'h45)? 32'h9d4d47cb
	         : (byte_in == 8'h46)? 32'h18c49f60
	         : (byte_in == 8'h47)? 32'hba598df7
	         : (byte_in == 8'h48)? 32'h5f35acae
	         : (byte_in == 8'h49)? 32'hfda8be39
	         : (byte_in == 8'h4a)? 32'h78216692
	         : (byte_in == 8'h4b)? 32'hdabc7405
	         : (byte_in == 8'h4c)? 32'hdff77a21
	         : (byte_in == 8'h4d)? 32'h7d6a68b6
	         : (byte_in == 8'h4e)? 32'hf8e3b01d
	         : (byte_in == 8'h4f)? 32'h5a7ea28a
	         : (byte_in == 8'h50)? 32'hd5606668
	         : (byte_in == 8'h51)? 32'h77fd74ff
	         : (byte_in == 8'h52)? 32'hf274ac54
	         : (byte_in == 8'h53)? 32'h50e9bec3
	         : (byte_in == 8'h54)? 32'h55a2b0e7
	         : (byte_in == 8'h55)? 32'hf73fa270
	         : (byte_in == 8'h56)? 32'h72b67adb
	         : (byte_in == 8'h57)? 32'hd02b684c
	         : (byte_in == 8'h58)? 32'h35474915
	         : (byte_in == 8'h59)? 32'h97da5b82
	         : (byte_in == 8'h5a)? 32'h12538329
	         : (byte_in == 8'h5b)? 32'hb0ce91be
	         : (byte_in == 8'h5c)? 32'hb5859f9a
	         : (byte_in == 8'h5d)? 32'h17188d0d
	         : (byte_in == 8'h5e)? 32'h929155a6
	         : (byte_in == 8'h5f)? 32'h300c4731
	         : (byte_in == 8'h60)? 32'hbaa52e89
	         : (byte_in == 8'h61)? 32'h18383c1e
	         : (byte_in == 8'h62)? 32'h9db1e4b5
	         : (byte_in == 8'h63)? 32'h3f2cf622
	         : (byte_in == 8'h64)? 32'h3a67f806
	         : (byte_in == 8'h65)? 32'h98faea91
	         : (byte_in == 8'h66)? 32'h1d73323a
	         : (byte_in == 8'h67)? 32'hbfee20ad
	         : (byte_in == 8'h68)? 32'h5a8201f4
	         : (byte_in == 8'h69)? 32'hf81f1363
	         : (byte_in == 8'h6a)? 32'h7d96cbc8
	         : (byte_in == 8'h6b)? 32'hdf0bd95f
	         : (byte_in == 8'h6c)? 32'hda40d77b
	         : (byte_in == 8'h6d)? 32'h78ddc5ec
	         : (byte_in == 8'h6e)? 32'hfd541d47
	         : (byte_in == 8'h6f)? 32'h5fc90fd0
	         : (byte_in == 8'h70)? 32'hd0d7cb32
	         : (byte_in == 8'h71)? 32'h724ad9a5
	         : (byte_in == 8'h72)? 32'hf7c3010e
	         : (byte_in == 8'h73)? 32'h555e1399
	         : (byte_in == 8'h74)? 32'h50151dbd
	         : (byte_in == 8'h75)? 32'hf2880f2a
	         : (byte_in == 8'h76)? 32'h7701d781
	         : (byte_in == 8'h77)? 32'hd59cc516
	         : (byte_in == 8'h78)? 32'h30f0e44f
	         : (byte_in == 8'h79)? 32'h926df6d8
	         : (byte_in == 8'h7a)? 32'h17e42e73
	         : (byte_in == 8'h7b)? 32'hb5793ce4
	         : (byte_in == 8'h7c)? 32'hb03232c0
	         : (byte_in == 8'h7d)? 32'h12af2057
	         : (byte_in == 8'h7e)? 32'h9726f8fc
	         : (byte_in == 8'h7f)? 32'h35bbea6b
	         : (byte_in == 8'h80)? 32'hce97a914
	         : (byte_in == 8'h81)? 32'h6c0abb83
	         : (byte_in == 8'h82)? 32'he9836328
	         : (byte_in == 8'h83)? 32'h4b1e71bf
	         : (byte_in == 8'h84)? 32'h4e557f9b
	         : (byte_in == 8'h85)? 32'hecc86d0c
	         : (byte_in == 8'h86)? 32'h6941b5a7
	         : (byte_in == 8'h87)? 32'hcbdca730
	         : (byte_in == 8'h88)? 32'h2eb08669
	         : (byte_in == 8'h89)? 32'h8c2d94fe
	         : (byte_in == 8'h8a)? 32'h09a44c55
	         : (byte_in == 8'h8b)? 32'hab395ec2
	         : (byte_in == 8'h8c)? 32'hae7250e6
	         : (byte_in == 8'h8d)? 32'h0cef4271
	         : (byte_in == 8'h8e)? 32'h89669ada
	         : (byte_in == 8'h8f)? 32'h2bfb884d
	         : (byte_in == 8'h90)? 32'ha4e54caf
	         : (byte_in == 8'h91)? 32'h06785e38
	         : (byte_in == 8'h92)? 32'h83f18693
	         : (byte_in == 8'h93)? 32'h216c9404
	         : (byte_in == 8'h94)? 32'h24279a20
	         : (byte_in == 8'h95)? 32'h86ba88b7
	         : (byte_in == 8'h96)? 32'h0333501c
	         : (byte_in == 8'h97)? 32'ha1ae428b
	         : (byte_in == 8'h98)? 32'h44c263d2
	         : (byte_in == 8'h99)? 32'he65f7145
	         : (byte_in == 8'h9a)? 32'h63d6a9ee
	         : (byte_in == 8'h9b)? 32'hc14bbb79
	         : (byte_in == 8'h9c)? 32'hc400b55d
	         : (byte_in == 8'h9d)? 32'h669da7ca
	         : (byte_in == 8'h9e)? 32'he3147f61
	         : (byte_in == 8'h9f)? 32'h41896df6
	         : (byte_in == 8'ha0)? 32'hcb20044e
	         : (byte_in == 8'ha1)? 32'h69bd16d9
	         : (byte_in == 8'ha2)? 32'hec34ce72
	         : (byte_in == 8'ha3)? 32'h4ea9dce5
	         : (byte_in == 8'ha4)? 32'h4be2d2c1
	         : (byte_in == 8'ha5)? 32'he97fc056
	         : (byte_in == 8'ha6)? 32'h6cf618fd
	         : (byte_in == 8'ha7)? 32'hce6b0a6a
	         : (byte_in == 8'ha8)? 32'h2b072b33
	         : (byte_in == 8'ha9)? 32'h899a39a4
	         : (byte_in == 8'haa)? 32'h0c13e10f
	         : (byte_in == 8'hab)? 32'hae8ef398
	         : (byte_in == 8'hac)? 32'habc5fdbc
	         : (byte_in == 8'had)? 32'h0958ef2b
	         : (byte_in == 8'hae)? 32'h8cd13780
	         : (byte_in == 8'haf)? 32'h2e4c2517
	         : (byte_in == 8'hb0)? 32'ha152e1f5
	         : (byte_in == 8'hb1)? 32'h03cff362
	         : (byte_in == 8'hb2)? 32'h86462bc9
	         : (byte_in == 8'hb3)? 32'h24db395e
	         : (byte_in == 8'hb4)? 32'h2190377a
	         : (byte_in == 8'hb5)? 32'h830d25ed
	         : (byte_in == 8'hb6)? 32'h0684fd46
	         : (byte_in == 8'hb7)? 32'ha419efd1
	         : (byte_in == 8'hb8)? 32'h4175ce88
	         : (byte_in == 8'hb9)? 32'he3e8dc1f
	         : (byte_in == 8'hba)? 32'h666104b4
	         : (byte_in == 8'hbb)? 32'hc4fc1623
	         : (byte_in == 8'hbc)? 32'hc1b71807
	         : (byte_in == 8'hbd)? 32'h632a0a90
	         : (byte_in == 8'hbe)? 32'he6a3d23b
	         : (byte_in == 8'hbf)? 32'h443ec0ac
	         : (byte_in == 8'hc0)? 32'h71852ac7
	         : (byte_in == 8'hc1)? 32'hd3183850
	         : (byte_in == 8'hc2)? 32'h5691e0fb
	         : (byte_in == 8'hc3)? 32'hf40cf26c
	         : (byte_in == 8'hc4)? 32'hf147fc48
	         : (byte_in == 8'hc5)? 32'h53daeedf
	         : (byte_in == 8'hc6)? 32'hd6533674
	         : (byte_in == 8'hc7)? 32'h74ce24e3
	         : (byte_in == 8'hc8)? 32'h91a205ba
	         : (byte_in == 8'hc9)? 32'h333f172d
	         : (byte_in == 8'hca)? 32'hb6b6cf86
	         : (byte_in == 8'hcb)? 32'h142bdd11
	         : (byte_in == 8'hcc)? 32'h1160d335
	         : (byte_in == 8'hcd)? 32'hb3fdc1a2
	         : (byte_in == 8'hce)? 32'h36741909
	         : (byte_in == 8'hcf)? 32'h94e90b9e
	         : (byte_in == 8'hd0)? 32'h1bf7cf7c
	         : (byte_in == 8'hd1)? 32'hb96addeb
	         : (byte_in == 8'hd2)? 32'h3ce30540
	         : (byte_in == 8'hd3)? 32'h9e7e17d7
	         : (byte_in == 8'hd4)? 32'h9b3519f3
	         : (byte_in == 8'hd5)? 32'h39a80b64
	         : (byte_in == 8'hd6)? 32'hbc21d3cf
	         : (byte_in == 8'hd7)? 32'h1ebcc158
	         : (byte_in == 8'hd8)? 32'hfbd0e001
	         : (byte_in == 8'hd9)? 32'h594df296
	         : (byte_in == 8'hda)? 32'hdcc42a3d
	         : (byte_in == 8'hdb)? 32'h7e5938aa
	         : (byte_in == 8'hdc)? 32'h7b12368e
	         : (byte_in == 8'hdd)? 32'hd98f2419
	         : (byte_in == 8'hde)? 32'h5c06fcb2
	         : (byte_in == 8'hdf)? 32'hfe9bee25
	         : (byte_in == 8'he0)? 32'h7432879d
	         : (byte_in == 8'he1)? 32'hd6af950a
	         : (byte_in == 8'he2)? 32'h53264da1
	         : (byte_in == 8'he3)? 32'hf1bb5f36
	         : (byte_in == 8'he4)? 32'hf4f05112
	         : (byte_in == 8'he5)? 32'h566d4385
	         : (byte_in == 8'he6)? 32'hd3e49b2e
	         : (byte_in == 8'he7)? 32'h717989b9
	         : (byte_in == 8'he8)? 32'h9415a8e0
	         : (byte_in == 8'he9)? 32'h3688ba77
	         : (byte_in == 8'hea)? 32'hb30162dc
	         : (byte_in == 8'heb)? 32'h119c704b
	         : (byte_in == 8'hec)? 32'h14d77e6f
	         : (byte_in == 8'hed)? 32'hb64a6cf8
	         : (byte_in == 8'hee)? 32'h33c3b453
	         : (byte_in == 8'hef)? 32'h915ea6c4
	         : (byte_in == 8'hf0)? 32'h1e406226
	         : (byte_in == 8'hf1)? 32'hbcdd70b1
	         : (byte_in == 8'hf2)? 32'h3954a81a
	         : (byte_in == 8'hf3)? 32'h9bc9ba8d
	         : (byte_in == 8'hf4)? 32'h9e82b4a9
	         : (byte_in == 8'hf5)? 32'h3c1fa63e
	         : (byte_in == 8'hf6)? 32'hb9967e95
	         : (byte_in == 8'hf7)? 32'h1b0b6c02
	         : (byte_in == 8'hf8)? 32'hfe674d5b
	         : (byte_in == 8'hf9)? 32'h5cfa5fcc
	         : (byte_in == 8'hfa)? 32'hd9738767
	         : (byte_in == 8'hfb)? 32'h7bee95f0
	         : (byte_in == 8'hfc)? 32'h7ea59bd4
	         : (byte_in == 8'hfd)? 32'hdc388943
	         : (byte_in == 8'hfe)? 32'h59b151e8
	         :                     32'hfb2c437f;

endmodule
//}}}

module TABLE27(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'hbbdcf407
	         : (byte_in == 8'h02)? 32'h3321e92c
	         : (byte_in == 8'h03)? 32'h88fd1d2b
	         : (byte_in == 8'h04)? 32'h77b9e80f
	         : (byte_in == 8'h05)? 32'hcc651c08
	         : (byte_in == 8'h06)? 32'h44980123
	         : (byte_in == 8'h07)? 32'hff44f524
	         : (byte_in == 8'h08)? 32'h6643d258
	         : (byte_in == 8'h09)? 32'hdd9f265f
	         : (byte_in == 8'h0a)? 32'h55623b74
	         : (byte_in == 8'h0b)? 32'heebecf73
	         : (byte_in == 8'h0c)? 32'h11fa3a57
	         : (byte_in == 8'h0d)? 32'haa26ce50
	         : (byte_in == 8'h0e)? 32'h22dbd37b
	         : (byte_in == 8'h0f)? 32'h9907277c
	         : (byte_in == 8'h10)? 32'h848598ba
	         : (byte_in == 8'h11)? 32'h3f596cbd
	         : (byte_in == 8'h12)? 32'hb7a47196
	         : (byte_in == 8'h13)? 32'h0c788591
	         : (byte_in == 8'h14)? 32'hf33c70b5
	         : (byte_in == 8'h15)? 32'h48e084b2
	         : (byte_in == 8'h16)? 32'hc01d9999
	         : (byte_in == 8'h17)? 32'h7bc16d9e
	         : (byte_in == 8'h18)? 32'he2c64ae2
	         : (byte_in == 8'h19)? 32'h591abee5
	         : (byte_in == 8'h1a)? 32'hd1e7a3ce
	         : (byte_in == 8'h1b)? 32'h6a3b57c9
	         : (byte_in == 8'h1c)? 32'h957fa2ed
	         : (byte_in == 8'h1d)? 32'h2ea356ea
	         : (byte_in == 8'h1e)? 32'ha65e4bc1
	         : (byte_in == 8'h1f)? 32'h1d82bfc6
	         : (byte_in == 8'h20)? 32'h097f5711
	         : (byte_in == 8'h21)? 32'hb2a3a316
	         : (byte_in == 8'h22)? 32'h3a5ebe3d
	         : (byte_in == 8'h23)? 32'h81824a3a
	         : (byte_in == 8'h24)? 32'h7ec6bf1e
	         : (byte_in == 8'h25)? 32'hc51a4b19
	         : (byte_in == 8'h26)? 32'h4de75632
	         : (byte_in == 8'h27)? 32'hf63ba235
	         : (byte_in == 8'h28)? 32'h6f3c8549
	         : (byte_in == 8'h29)? 32'hd4e0714e
	         : (byte_in == 8'h2a)? 32'h5c1d6c65
	         : (byte_in == 8'h2b)? 32'he7c19862
	         : (byte_in == 8'h2c)? 32'h18856d46
	         : (byte_in == 8'h2d)? 32'ha3599941
	         : (byte_in == 8'h2e)? 32'h2ba4846a
	         : (byte_in == 8'h2f)? 32'h9078706d
	         : (byte_in == 8'h30)? 32'h8dfacfab
	         : (byte_in == 8'h31)? 32'h36263bac
	         : (byte_in == 8'h32)? 32'hbedb2687
	         : (byte_in == 8'h33)? 32'h0507d280
	         : (byte_in == 8'h34)? 32'hfa4327a4
	         : (byte_in == 8'h35)? 32'h419fd3a3
	         : (byte_in == 8'h36)? 32'hc962ce88
	         : (byte_in == 8'h37)? 32'h72be3a8f
	         : (byte_in == 8'h38)? 32'hebb91df3
	         : (byte_in == 8'h39)? 32'h5065e9f4
	         : (byte_in == 8'h3a)? 32'hd898f4df
	         : (byte_in == 8'h3b)? 32'h634400d8
	         : (byte_in == 8'h3c)? 32'h9c00f5fc
	         : (byte_in == 8'h3d)? 32'h27dc01fb
	         : (byte_in == 8'h3e)? 32'haf211cd0
	         : (byte_in == 8'h3f)? 32'h14fde8d7
	         : (byte_in == 8'h40)? 32'h62fc79d0
	         : (byte_in == 8'h41)? 32'hd9208dd7
	         : (byte_in == 8'h42)? 32'h51dd90fc
	         : (byte_in == 8'h43)? 32'hea0164fb
	         : (byte_in == 8'h44)? 32'h154591df
	         : (byte_in == 8'h45)? 32'hae9965d8
	         : (byte_in == 8'h46)? 32'h266478f3
	         : (byte_in == 8'h47)? 32'h9db88cf4
	         : (byte_in == 8'h48)? 32'h04bfab88
	         : (byte_in == 8'h49)? 32'hbf635f8f
	         : (byte_in == 8'h4a)? 32'h379e42a4
	         : (byte_in == 8'h4b)? 32'h8c42b6a3
	         : (byte_in == 8'h4c)? 32'h73064387
	         : (byte_in == 8'h4d)? 32'hc8dab780
	         : (byte_in == 8'h4e)? 32'h4027aaab
	         : (byte_in == 8'h4f)? 32'hfbfb5eac
	         : (byte_in == 8'h50)? 32'he679e16a
	         : (byte_in == 8'h51)? 32'h5da5156d
	         : (byte_in == 8'h52)? 32'hd5580846
	         : (byte_in == 8'h53)? 32'h6e84fc41
	         : (byte_in == 8'h54)? 32'h91c00965
	         : (byte_in == 8'h55)? 32'h2a1cfd62
	         : (byte_in == 8'h56)? 32'ha2e1e049
	         : (byte_in == 8'h57)? 32'h193d144e
	         : (byte_in == 8'h58)? 32'h803a3332
	         : (byte_in == 8'h59)? 32'h3be6c735
	         : (byte_in == 8'h5a)? 32'hb31bda1e
	         : (byte_in == 8'h5b)? 32'h08c72e19
	         : (byte_in == 8'h5c)? 32'hf783db3d
	         : (byte_in == 8'h5d)? 32'h4c5f2f3a
	         : (byte_in == 8'h5e)? 32'hc4a23211
	         : (byte_in == 8'h5f)? 32'h7f7ec616
	         : (byte_in == 8'h60)? 32'h6b832ec1
	         : (byte_in == 8'h61)? 32'hd05fdac6
	         : (byte_in == 8'h62)? 32'h58a2c7ed
	         : (byte_in == 8'h63)? 32'he37e33ea
	         : (byte_in == 8'h64)? 32'h1c3ac6ce
	         : (byte_in == 8'h65)? 32'ha7e632c9
	         : (byte_in == 8'h66)? 32'h2f1b2fe2
	         : (byte_in == 8'h67)? 32'h94c7dbe5
	         : (byte_in == 8'h68)? 32'h0dc0fc99
	         : (byte_in == 8'h69)? 32'hb61c089e
	         : (byte_in == 8'h6a)? 32'h3ee115b5
	         : (byte_in == 8'h6b)? 32'h853de1b2
	         : (byte_in == 8'h6c)? 32'h7a791496
	         : (byte_in == 8'h6d)? 32'hc1a5e091
	         : (byte_in == 8'h6e)? 32'h4958fdba
	         : (byte_in == 8'h6f)? 32'hf28409bd
	         : (byte_in == 8'h70)? 32'hef06b67b
	         : (byte_in == 8'h71)? 32'h54da427c
	         : (byte_in == 8'h72)? 32'hdc275f57
	         : (byte_in == 8'h73)? 32'h67fbab50
	         : (byte_in == 8'h74)? 32'h98bf5e74
	         : (byte_in == 8'h75)? 32'h2363aa73
	         : (byte_in == 8'h76)? 32'hab9eb758
	         : (byte_in == 8'h77)? 32'h1042435f
	         : (byte_in == 8'h78)? 32'h89456423
	         : (byte_in == 8'h79)? 32'h32999024
	         : (byte_in == 8'h7a)? 32'hba648d0f
	         : (byte_in == 8'h7b)? 32'h01b87908
	         : (byte_in == 8'h7c)? 32'hfefc8c2c
	         : (byte_in == 8'h7d)? 32'h4520782b
	         : (byte_in == 8'h7e)? 32'hcddd6500
	         : (byte_in == 8'h7f)? 32'h76019107
	         : (byte_in == 8'h80)? 32'hd7075d82
	         : (byte_in == 8'h81)? 32'h6cdba985
	         : (byte_in == 8'h82)? 32'he426b4ae
	         : (byte_in == 8'h83)? 32'h5ffa40a9
	         : (byte_in == 8'h84)? 32'ha0beb58d
	         : (byte_in == 8'h85)? 32'h1b62418a
	         : (byte_in == 8'h86)? 32'h939f5ca1
	         : (byte_in == 8'h87)? 32'h2843a8a6
	         : (byte_in == 8'h88)? 32'hb1448fda
	         : (byte_in == 8'h89)? 32'h0a987bdd
	         : (byte_in == 8'h8a)? 32'h826566f6
	         : (byte_in == 8'h8b)? 32'h39b992f1
	         : (byte_in == 8'h8c)? 32'hc6fd67d5
	         : (byte_in == 8'h8d)? 32'h7d2193d2
	         : (byte_in == 8'h8e)? 32'hf5dc8ef9
	         : (byte_in == 8'h8f)? 32'h4e007afe
	         : (byte_in == 8'h90)? 32'h5382c538
	         : (byte_in == 8'h91)? 32'he85e313f
	         : (byte_in == 8'h92)? 32'h60a32c14
	         : (byte_in == 8'h93)? 32'hdb7fd813
	         : (byte_in == 8'h94)? 32'h243b2d37
	         : (byte_in == 8'h95)? 32'h9fe7d930
	         : (byte_in == 8'h96)? 32'h171ac41b
	         : (byte_in == 8'h97)? 32'hacc6301c
	         : (byte_in == 8'h98)? 32'h35c11760
	         : (byte_in == 8'h99)? 32'h8e1de367
	         : (byte_in == 8'h9a)? 32'h06e0fe4c
	         : (byte_in == 8'h9b)? 32'hbd3c0a4b
	         : (byte_in == 8'h9c)? 32'h4278ff6f
	         : (byte_in == 8'h9d)? 32'hf9a40b68
	         : (byte_in == 8'h9e)? 32'h71591643
	         : (byte_in == 8'h9f)? 32'hca85e244
	         : (byte_in == 8'ha0)? 32'hde780a93
	         : (byte_in == 8'ha1)? 32'h65a4fe94
	         : (byte_in == 8'ha2)? 32'hed59e3bf
	         : (byte_in == 8'ha3)? 32'h568517b8
	         : (byte_in == 8'ha4)? 32'ha9c1e29c
	         : (byte_in == 8'ha5)? 32'h121d169b
	         : (byte_in == 8'ha6)? 32'h9ae00bb0
	         : (byte_in == 8'ha7)? 32'h213cffb7
	         : (byte_in == 8'ha8)? 32'hb83bd8cb
	         : (byte_in == 8'ha9)? 32'h03e72ccc
	         : (byte_in == 8'haa)? 32'h8b1a31e7
	         : (byte_in == 8'hab)? 32'h30c6c5e0
	         : (byte_in == 8'hac)? 32'hcf8230c4
	         : (byte_in == 8'had)? 32'h745ec4c3
	         : (byte_in == 8'hae)? 32'hfca3d9e8
	         : (byte_in == 8'haf)? 32'h477f2def
	         : (byte_in == 8'hb0)? 32'h5afd9229
	         : (byte_in == 8'hb1)? 32'he121662e
	         : (byte_in == 8'hb2)? 32'h69dc7b05
	         : (byte_in == 8'hb3)? 32'hd2008f02
	         : (byte_in == 8'hb4)? 32'h2d447a26
	         : (byte_in == 8'hb5)? 32'h96988e21
	         : (byte_in == 8'hb6)? 32'h1e65930a
	         : (byte_in == 8'hb7)? 32'ha5b9670d
	         : (byte_in == 8'hb8)? 32'h3cbe4071
	         : (byte_in == 8'hb9)? 32'h8762b476
	         : (byte_in == 8'hba)? 32'h0f9fa95d
	         : (byte_in == 8'hbb)? 32'hb4435d5a
	         : (byte_in == 8'hbc)? 32'h4b07a87e
	         : (byte_in == 8'hbd)? 32'hf0db5c79
	         : (byte_in == 8'hbe)? 32'h78264152
	         : (byte_in == 8'hbf)? 32'hc3fab555
	         : (byte_in == 8'hc0)? 32'hb5fb2452
	         : (byte_in == 8'hc1)? 32'h0e27d055
	         : (byte_in == 8'hc2)? 32'h86dacd7e
	         : (byte_in == 8'hc3)? 32'h3d063979
	         : (byte_in == 8'hc4)? 32'hc242cc5d
	         : (byte_in == 8'hc5)? 32'h799e385a
	         : (byte_in == 8'hc6)? 32'hf1632571
	         : (byte_in == 8'hc7)? 32'h4abfd176
	         : (byte_in == 8'hc8)? 32'hd3b8f60a
	         : (byte_in == 8'hc9)? 32'h6864020d
	         : (byte_in == 8'hca)? 32'he0991f26
	         : (byte_in == 8'hcb)? 32'h5b45eb21
	         : (byte_in == 8'hcc)? 32'ha4011e05
	         : (byte_in == 8'hcd)? 32'h1fddea02
	         : (byte_in == 8'hce)? 32'h9720f729
	         : (byte_in == 8'hcf)? 32'h2cfc032e
	         : (byte_in == 8'hd0)? 32'h317ebce8
	         : (byte_in == 8'hd1)? 32'h8aa248ef
	         : (byte_in == 8'hd2)? 32'h025f55c4
	         : (byte_in == 8'hd3)? 32'hb983a1c3
	         : (byte_in == 8'hd4)? 32'h46c754e7
	         : (byte_in == 8'hd5)? 32'hfd1ba0e0
	         : (byte_in == 8'hd6)? 32'h75e6bdcb
	         : (byte_in == 8'hd7)? 32'hce3a49cc
	         : (byte_in == 8'hd8)? 32'h573d6eb0
	         : (byte_in == 8'hd9)? 32'hece19ab7
	         : (byte_in == 8'hda)? 32'h641c879c
	         : (byte_in == 8'hdb)? 32'hdfc0739b
	         : (byte_in == 8'hdc)? 32'h208486bf
	         : (byte_in == 8'hdd)? 32'h9b5872b8
	         : (byte_in == 8'hde)? 32'h13a56f93
	         : (byte_in == 8'hdf)? 32'ha8799b94
	         : (byte_in == 8'he0)? 32'hbc847343
	         : (byte_in == 8'he1)? 32'h07588744
	         : (byte_in == 8'he2)? 32'h8fa59a6f
	         : (byte_in == 8'he3)? 32'h34796e68
	         : (byte_in == 8'he4)? 32'hcb3d9b4c
	         : (byte_in == 8'he5)? 32'h70e16f4b
	         : (byte_in == 8'he6)? 32'hf81c7260
	         : (byte_in == 8'he7)? 32'h43c08667
	         : (byte_in == 8'he8)? 32'hdac7a11b
	         : (byte_in == 8'he9)? 32'h611b551c
	         : (byte_in == 8'hea)? 32'he9e64837
	         : (byte_in == 8'heb)? 32'h523abc30
	         : (byte_in == 8'hec)? 32'had7e4914
	         : (byte_in == 8'hed)? 32'h16a2bd13
	         : (byte_in == 8'hee)? 32'h9e5fa038
	         : (byte_in == 8'hef)? 32'h2583543f
	         : (byte_in == 8'hf0)? 32'h3801ebf9
	         : (byte_in == 8'hf1)? 32'h83dd1ffe
	         : (byte_in == 8'hf2)? 32'h0b2002d5
	         : (byte_in == 8'hf3)? 32'hb0fcf6d2
	         : (byte_in == 8'hf4)? 32'h4fb803f6
	         : (byte_in == 8'hf5)? 32'hf464f7f1
	         : (byte_in == 8'hf6)? 32'h7c99eada
	         : (byte_in == 8'hf7)? 32'hc7451edd
	         : (byte_in == 8'hf8)? 32'h5e4239a1
	         : (byte_in == 8'hf9)? 32'he59ecda6
	         : (byte_in == 8'hfa)? 32'h6d63d08d
	         : (byte_in == 8'hfb)? 32'hd6bf248a
	         : (byte_in == 8'hfc)? 32'h29fbd1ae
	         : (byte_in == 8'hfd)? 32'h922725a9
	         : (byte_in == 8'hfe)? 32'h1ada3882
	         :                     32'ha106cc85;

endmodule
//}}}

module TABLE28(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h539cbdbf
	         : (byte_in == 8'h02)? 32'he6387b84
	         : (byte_in == 8'h03)? 32'hb5a4c63b
	         : (byte_in == 8'h04)? 32'h1298bd46
	         : (byte_in == 8'h05)? 32'h410400f9
	         : (byte_in == 8'h06)? 32'hf4a0c6c2
	         : (byte_in == 8'h07)? 32'ha73c7b7d
	         : (byte_in == 8'h08)? 32'h9fed4ab7
	         : (byte_in == 8'h09)? 32'hcc71f708
	         : (byte_in == 8'h0a)? 32'h79d53133
	         : (byte_in == 8'h0b)? 32'h2a498c8c
	         : (byte_in == 8'h0c)? 32'h8d75f7f1
	         : (byte_in == 8'h0d)? 32'hdee94a4e
	         : (byte_in == 8'h0e)? 32'h6b4d8c75
	         : (byte_in == 8'h0f)? 32'h38d131ca
	         : (byte_in == 8'h10)? 32'h76acc733
	         : (byte_in == 8'h11)? 32'h25307a8c
	         : (byte_in == 8'h12)? 32'h9094bcb7
	         : (byte_in == 8'h13)? 32'hc3080108
	         : (byte_in == 8'h14)? 32'h64347a75
	         : (byte_in == 8'h15)? 32'h37a8c7ca
	         : (byte_in == 8'h16)? 32'h820c01f1
	         : (byte_in == 8'h17)? 32'hd190bc4e
	         : (byte_in == 8'h18)? 32'he9418d84
	         : (byte_in == 8'h19)? 32'hbadd303b
	         : (byte_in == 8'h1a)? 32'h0f79f600
	         : (byte_in == 8'h1b)? 32'h5ce54bbf
	         : (byte_in == 8'h1c)? 32'hfbd930c2
	         : (byte_in == 8'h1d)? 32'ha8458d7d
	         : (byte_in == 8'h1e)? 32'h1de14b46
	         : (byte_in == 8'h1f)? 32'h4e7df6f9
	         : (byte_in == 8'h20)? 32'hd9e6eee9
	         : (byte_in == 8'h21)? 32'h8a7a5356
	         : (byte_in == 8'h22)? 32'h3fde956d
	         : (byte_in == 8'h23)? 32'h6c4228d2
	         : (byte_in == 8'h24)? 32'hcb7e53af
	         : (byte_in == 8'h25)? 32'h98e2ee10
	         : (byte_in == 8'h26)? 32'h2d46282b
	         : (byte_in == 8'h27)? 32'h7eda9594
	         : (byte_in == 8'h28)? 32'h460ba45e
	         : (byte_in == 8'h29)? 32'h159719e1
	         : (byte_in == 8'h2a)? 32'ha033dfda
	         : (byte_in == 8'h2b)? 32'hf3af6265
	         : (byte_in == 8'h2c)? 32'h54931918
	         : (byte_in == 8'h2d)? 32'h070fa4a7
	         : (byte_in == 8'h2e)? 32'hb2ab629c
	         : (byte_in == 8'h2f)? 32'he137df23
	         : (byte_in == 8'h30)? 32'haf4a29da
	         : (byte_in == 8'h31)? 32'hfcd69465
	         : (byte_in == 8'h32)? 32'h4972525e
	         : (byte_in == 8'h33)? 32'h1aeeefe1
	         : (byte_in == 8'h34)? 32'hbdd2949c
	         : (byte_in == 8'h35)? 32'hee4e2923
	         : (byte_in == 8'h36)? 32'h5beaef18
	         : (byte_in == 8'h37)? 32'h087652a7
	         : (byte_in == 8'h38)? 32'h30a7636d
	         : (byte_in == 8'h39)? 32'h633bded2
	         : (byte_in == 8'h3a)? 32'hd69f18e9
	         : (byte_in == 8'h3b)? 32'h8503a556
	         : (byte_in == 8'h3c)? 32'h223fde2b
	         : (byte_in == 8'h3d)? 32'h71a36394
	         : (byte_in == 8'h3e)? 32'hc407a5af
	         : (byte_in == 8'h3f)? 32'h979b1810
	         : (byte_in == 8'h40)? 32'h58f8485f
	         : (byte_in == 8'h41)? 32'h0b64f5e0
	         : (byte_in == 8'h42)? 32'hbec033db
	         : (byte_in == 8'h43)? 32'hed5c8e64
	         : (byte_in == 8'h44)? 32'h4a60f519
	         : (byte_in == 8'h45)? 32'h19fc48a6
	         : (byte_in == 8'h46)? 32'hac588e9d
	         : (byte_in == 8'h47)? 32'hffc43322
	         : (byte_in == 8'h48)? 32'hc71502e8
	         : (byte_in == 8'h49)? 32'h9489bf57
	         : (byte_in == 8'h4a)? 32'h212d796c
	         : (byte_in == 8'h4b)? 32'h72b1c4d3
	         : (byte_in == 8'h4c)? 32'hd58dbfae
	         : (byte_in == 8'h4d)? 32'h86110211
	         : (byte_in == 8'h4e)? 32'h33b5c42a
	         : (byte_in == 8'h4f)? 32'h60297995
	         : (byte_in == 8'h50)? 32'h2e548f6c
	         : (byte_in == 8'h51)? 32'h7dc832d3
	         : (byte_in == 8'h52)? 32'hc86cf4e8
	         : (byte_in == 8'h53)? 32'h9bf04957
	         : (byte_in == 8'h54)? 32'h3ccc322a
	         : (byte_in == 8'h55)? 32'h6f508f95
	         : (byte_in == 8'h56)? 32'hdaf449ae
	         : (byte_in == 8'h57)? 32'h8968f411
	         : (byte_in == 8'h58)? 32'hb1b9c5db
	         : (byte_in == 8'h59)? 32'he2257864
	         : (byte_in == 8'h5a)? 32'h5781be5f
	         : (byte_in == 8'h5b)? 32'h041d03e0
	         : (byte_in == 8'h5c)? 32'ha321789d
	         : (byte_in == 8'h5d)? 32'hf0bdc522
	         : (byte_in == 8'h5e)? 32'h45190319
	         : (byte_in == 8'h5f)? 32'h1685bea6
	         : (byte_in == 8'h60)? 32'h811ea6b6
	         : (byte_in == 8'h61)? 32'hd2821b09
	         : (byte_in == 8'h62)? 32'h6726dd32
	         : (byte_in == 8'h63)? 32'h34ba608d
	         : (byte_in == 8'h64)? 32'h93861bf0
	         : (byte_in == 8'h65)? 32'hc01aa64f
	         : (byte_in == 8'h66)? 32'h75be6074
	         : (byte_in == 8'h67)? 32'h2622ddcb
	         : (byte_in == 8'h68)? 32'h1ef3ec01
	         : (byte_in == 8'h69)? 32'h4d6f51be
	         : (byte_in == 8'h6a)? 32'hf8cb9785
	         : (byte_in == 8'h6b)? 32'hab572a3a
	         : (byte_in == 8'h6c)? 32'h0c6b5147
	         : (byte_in == 8'h6d)? 32'h5ff7ecf8
	         : (byte_in == 8'h6e)? 32'hea532ac3
	         : (byte_in == 8'h6f)? 32'hb9cf977c
	         : (byte_in == 8'h70)? 32'hf7b26185
	         : (byte_in == 8'h71)? 32'ha42edc3a
	         : (byte_in == 8'h72)? 32'h118a1a01
	         : (byte_in == 8'h73)? 32'h4216a7be
	         : (byte_in == 8'h74)? 32'he52adcc3
	         : (byte_in == 8'h75)? 32'hb6b6617c
	         : (byte_in == 8'h76)? 32'h0312a747
	         : (byte_in == 8'h77)? 32'h508e1af8
	         : (byte_in == 8'h78)? 32'h685f2b32
	         : (byte_in == 8'h79)? 32'h3bc3968d
	         : (byte_in == 8'h7a)? 32'h8e6750b6
	         : (byte_in == 8'h7b)? 32'hddfbed09
	         : (byte_in == 8'h7c)? 32'h7ac79674
	         : (byte_in == 8'h7d)? 32'h295b2bcb
	         : (byte_in == 8'h7e)? 32'h9cffedf0
	         : (byte_in == 8'h7f)? 32'hcf63504f
	         : (byte_in == 8'h80)? 32'he051606e
	         : (byte_in == 8'h81)? 32'hb3cdddd1
	         : (byte_in == 8'h82)? 32'h06691bea
	         : (byte_in == 8'h83)? 32'h55f5a655
	         : (byte_in == 8'h84)? 32'hf2c9dd28
	         : (byte_in == 8'h85)? 32'ha1556097
	         : (byte_in == 8'h86)? 32'h14f1a6ac
	         : (byte_in == 8'h87)? 32'h476d1b13
	         : (byte_in == 8'h88)? 32'h7fbc2ad9
	         : (byte_in == 8'h89)? 32'h2c209766
	         : (byte_in == 8'h8a)? 32'h9984515d
	         : (byte_in == 8'h8b)? 32'hca18ece2
	         : (byte_in == 8'h8c)? 32'h6d24979f
	         : (byte_in == 8'h8d)? 32'h3eb82a20
	         : (byte_in == 8'h8e)? 32'h8b1cec1b
	         : (byte_in == 8'h8f)? 32'hd88051a4
	         : (byte_in == 8'h90)? 32'h96fda75d
	         : (byte_in == 8'h91)? 32'hc5611ae2
	         : (byte_in == 8'h92)? 32'h70c5dcd9
	         : (byte_in == 8'h93)? 32'h23596166
	         : (byte_in == 8'h94)? 32'h84651a1b
	         : (byte_in == 8'h95)? 32'hd7f9a7a4
	         : (byte_in == 8'h96)? 32'h625d619f
	         : (byte_in == 8'h97)? 32'h31c1dc20
	         : (byte_in == 8'h98)? 32'h0910edea
	         : (byte_in == 8'h99)? 32'h5a8c5055
	         : (byte_in == 8'h9a)? 32'hef28966e
	         : (byte_in == 8'h9b)? 32'hbcb42bd1
	         : (byte_in == 8'h9c)? 32'h1b8850ac
	         : (byte_in == 8'h9d)? 32'h4814ed13
	         : (byte_in == 8'h9e)? 32'hfdb02b28
	         : (byte_in == 8'h9f)? 32'hae2c9697
	         : (byte_in == 8'ha0)? 32'h39b78e87
	         : (byte_in == 8'ha1)? 32'h6a2b3338
	         : (byte_in == 8'ha2)? 32'hdf8ff503
	         : (byte_in == 8'ha3)? 32'h8c1348bc
	         : (byte_in == 8'ha4)? 32'h2b2f33c1
	         : (byte_in == 8'ha5)? 32'h78b38e7e
	         : (byte_in == 8'ha6)? 32'hcd174845
	         : (byte_in == 8'ha7)? 32'h9e8bf5fa
	         : (byte_in == 8'ha8)? 32'ha65ac430
	         : (byte_in == 8'ha9)? 32'hf5c6798f
	         : (byte_in == 8'haa)? 32'h4062bfb4
	         : (byte_in == 8'hab)? 32'h13fe020b
	         : (byte_in == 8'hac)? 32'hb4c27976
	         : (byte_in == 8'had)? 32'he75ec4c9
	         : (byte_in == 8'hae)? 32'h52fa02f2
	         : (byte_in == 8'haf)? 32'h0166bf4d
	         : (byte_in == 8'hb0)? 32'h4f1b49b4
	         : (byte_in == 8'hb1)? 32'h1c87f40b
	         : (byte_in == 8'hb2)? 32'ha9233230
	         : (byte_in == 8'hb3)? 32'hfabf8f8f
	         : (byte_in == 8'hb4)? 32'h5d83f4f2
	         : (byte_in == 8'hb5)? 32'h0e1f494d
	         : (byte_in == 8'hb6)? 32'hbbbb8f76
	         : (byte_in == 8'hb7)? 32'he82732c9
	         : (byte_in == 8'hb8)? 32'hd0f60303
	         : (byte_in == 8'hb9)? 32'h836abebc
	         : (byte_in == 8'hba)? 32'h36ce7887
	         : (byte_in == 8'hbb)? 32'h6552c538
	         : (byte_in == 8'hbc)? 32'hc26ebe45
	         : (byte_in == 8'hbd)? 32'h91f203fa
	         : (byte_in == 8'hbe)? 32'h2456c5c1
	         : (byte_in == 8'hbf)? 32'h77ca787e
	         : (byte_in == 8'hc0)? 32'hb8a92831
	         : (byte_in == 8'hc1)? 32'heb35958e
	         : (byte_in == 8'hc2)? 32'h5e9153b5
	         : (byte_in == 8'hc3)? 32'h0d0dee0a
	         : (byte_in == 8'hc4)? 32'haa319577
	         : (byte_in == 8'hc5)? 32'hf9ad28c8
	         : (byte_in == 8'hc6)? 32'h4c09eef3
	         : (byte_in == 8'hc7)? 32'h1f95534c
	         : (byte_in == 8'hc8)? 32'h27446286
	         : (byte_in == 8'hc9)? 32'h74d8df39
	         : (byte_in == 8'hca)? 32'hc17c1902
	         : (byte_in == 8'hcb)? 32'h92e0a4bd
	         : (byte_in == 8'hcc)? 32'h35dcdfc0
	         : (byte_in == 8'hcd)? 32'h6640627f
	         : (byte_in == 8'hce)? 32'hd3e4a444
	         : (byte_in == 8'hcf)? 32'h807819fb
	         : (byte_in == 8'hd0)? 32'hce05ef02
	         : (byte_in == 8'hd1)? 32'h9d9952bd
	         : (byte_in == 8'hd2)? 32'h283d9486
	         : (byte_in == 8'hd3)? 32'h7ba12939
	         : (byte_in == 8'hd4)? 32'hdc9d5244
	         : (byte_in == 8'hd5)? 32'h8f01effb
	         : (byte_in == 8'hd6)? 32'h3aa529c0
	         : (byte_in == 8'hd7)? 32'h6939947f
	         : (byte_in == 8'hd8)? 32'h51e8a5b5
	         : (byte_in == 8'hd9)? 32'h0274180a
	         : (byte_in == 8'hda)? 32'hb7d0de31
	         : (byte_in == 8'hdb)? 32'he44c638e
	         : (byte_in == 8'hdc)? 32'h437018f3
	         : (byte_in == 8'hdd)? 32'h10eca54c
	         : (byte_in == 8'hde)? 32'ha5486377
	         : (byte_in == 8'hdf)? 32'hf6d4dec8
	         : (byte_in == 8'he0)? 32'h614fc6d8
	         : (byte_in == 8'he1)? 32'h32d37b67
	         : (byte_in == 8'he2)? 32'h8777bd5c
	         : (byte_in == 8'he3)? 32'hd4eb00e3
	         : (byte_in == 8'he4)? 32'h73d77b9e
	         : (byte_in == 8'he5)? 32'h204bc621
	         : (byte_in == 8'he6)? 32'h95ef001a
	         : (byte_in == 8'he7)? 32'hc673bda5
	         : (byte_in == 8'he8)? 32'hfea28c6f
	         : (byte_in == 8'he9)? 32'had3e31d0
	         : (byte_in == 8'hea)? 32'h189af7eb
	         : (byte_in == 8'heb)? 32'h4b064a54
	         : (byte_in == 8'hec)? 32'hec3a3129
	         : (byte_in == 8'hed)? 32'hbfa68c96
	         : (byte_in == 8'hee)? 32'h0a024aad
	         : (byte_in == 8'hef)? 32'h599ef712
	         : (byte_in == 8'hf0)? 32'h17e301eb
	         : (byte_in == 8'hf1)? 32'h447fbc54
	         : (byte_in == 8'hf2)? 32'hf1db7a6f
	         : (byte_in == 8'hf3)? 32'ha247c7d0
	         : (byte_in == 8'hf4)? 32'h057bbcad
	         : (byte_in == 8'hf5)? 32'h56e70112
	         : (byte_in == 8'hf6)? 32'he343c729
	         : (byte_in == 8'hf7)? 32'hb0df7a96
	         : (byte_in == 8'hf8)? 32'h880e4b5c
	         : (byte_in == 8'hf9)? 32'hdb92f6e3
	         : (byte_in == 8'hfa)? 32'h6e3630d8
	         : (byte_in == 8'hfb)? 32'h3daa8d67
	         : (byte_in == 8'hfc)? 32'h9a96f61a
	         : (byte_in == 8'hfd)? 32'hc90a4ba5
	         : (byte_in == 8'hfe)? 32'h7cae8d9e
	         :                     32'h2f323021;

endmodule
//}}}

module TABLE29(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'hb1f490bc
	         : (byte_in == 8'h02)? 32'hc0a3c0dd
	         : (byte_in == 8'h03)? 32'h71575061
	         : (byte_in == 8'h04)? 32'h63e92178
	         : (byte_in == 8'h05)? 32'hd21db1c4
	         : (byte_in == 8'h06)? 32'ha34ae1a5
	         : (byte_in == 8'h07)? 32'h12be7119
	         : (byte_in == 8'h08)? 32'h814681b8
	         : (byte_in == 8'h09)? 32'h30b21104
	         : (byte_in == 8'h0a)? 32'h41e54165
	         : (byte_in == 8'h0b)? 32'hf011d1d9
	         : (byte_in == 8'h0c)? 32'he2afa0c0
	         : (byte_in == 8'h0d)? 32'h535b307c
	         : (byte_in == 8'h0e)? 32'h220c601d
	         : (byte_in == 8'h0f)? 32'h93f8f0a1
	         : (byte_in == 8'h10)? 32'h727784cb
	         : (byte_in == 8'h11)? 32'hc3831477
	         : (byte_in == 8'h12)? 32'hb2d44416
	         : (byte_in == 8'h13)? 32'h0320d4aa
	         : (byte_in == 8'h14)? 32'h119ea5b3
	         : (byte_in == 8'h15)? 32'ha06a350f
	         : (byte_in == 8'h16)? 32'hd13d656e
	         : (byte_in == 8'h17)? 32'h60c9f5d2
	         : (byte_in == 8'h18)? 32'hf3310573
	         : (byte_in == 8'h19)? 32'h42c595cf
	         : (byte_in == 8'h1a)? 32'h3392c5ae
	         : (byte_in == 8'h1b)? 32'h82665512
	         : (byte_in == 8'h1c)? 32'h90d8240b
	         : (byte_in == 8'h1d)? 32'h212cb4b7
	         : (byte_in == 8'h1e)? 32'h507be4d6
	         : (byte_in == 8'h1f)? 32'he18f746a
	         : (byte_in == 8'h20)? 32'h5114bece
	         : (byte_in == 8'h21)? 32'he0e02e72
	         : (byte_in == 8'h22)? 32'h91b77e13
	         : (byte_in == 8'h23)? 32'h2043eeaf
	         : (byte_in == 8'h24)? 32'h32fd9fb6
	         : (byte_in == 8'h25)? 32'h83090f0a
	         : (byte_in == 8'h26)? 32'hf25e5f6b
	         : (byte_in == 8'h27)? 32'h43aacfd7
	         : (byte_in == 8'h28)? 32'hd0523f76
	         : (byte_in == 8'h29)? 32'h61a6afca
	         : (byte_in == 8'h2a)? 32'h10f1ffab
	         : (byte_in == 8'h2b)? 32'ha1056f17
	         : (byte_in == 8'h2c)? 32'hb3bb1e0e
	         : (byte_in == 8'h2d)? 32'h024f8eb2
	         : (byte_in == 8'h2e)? 32'h7318ded3
	         : (byte_in == 8'h2f)? 32'hc2ec4e6f
	         : (byte_in == 8'h30)? 32'h23633a05
	         : (byte_in == 8'h31)? 32'h9297aab9
	         : (byte_in == 8'h32)? 32'he3c0fad8
	         : (byte_in == 8'h33)? 32'h52346a64
	         : (byte_in == 8'h34)? 32'h408a1b7d
	         : (byte_in == 8'h35)? 32'hf17e8bc1
	         : (byte_in == 8'h36)? 32'h8029dba0
	         : (byte_in == 8'h37)? 32'h31dd4b1c
	         : (byte_in == 8'h38)? 32'ha225bbbd
	         : (byte_in == 8'h39)? 32'h13d12b01
	         : (byte_in == 8'h3a)? 32'h62867b60
	         : (byte_in == 8'h3b)? 32'hd372ebdc
	         : (byte_in == 8'h3c)? 32'hc1cc9ac5
	         : (byte_in == 8'h3d)? 32'h70380a79
	         : (byte_in == 8'h3e)? 32'h016f5a18
	         : (byte_in == 8'h3f)? 32'hb09bcaa4
	         : (byte_in == 8'h40)? 32'hb772b42b
	         : (byte_in == 8'h41)? 32'h06862497
	         : (byte_in == 8'h42)? 32'h77d174f6
	         : (byte_in == 8'h43)? 32'hc625e44a
	         : (byte_in == 8'h44)? 32'hd49b9553
	         : (byte_in == 8'h45)? 32'h656f05ef
	         : (byte_in == 8'h46)? 32'h1438558e
	         : (byte_in == 8'h47)? 32'ha5ccc532
	         : (byte_in == 8'h48)? 32'h36343593
	         : (byte_in == 8'h49)? 32'h87c0a52f
	         : (byte_in == 8'h4a)? 32'hf697f54e
	         : (byte_in == 8'h4b)? 32'h476365f2
	         : (byte_in == 8'h4c)? 32'h55dd14eb
	         : (byte_in == 8'h4d)? 32'he4298457
	         : (byte_in == 8'h4e)? 32'h957ed436
	         : (byte_in == 8'h4f)? 32'h248a448a
	         : (byte_in == 8'h50)? 32'hc50530e0
	         : (byte_in == 8'h51)? 32'h74f1a05c
	         : (byte_in == 8'h52)? 32'h05a6f03d
	         : (byte_in == 8'h53)? 32'hb4526081
	         : (byte_in == 8'h54)? 32'ha6ec1198
	         : (byte_in == 8'h55)? 32'h17188124
	         : (byte_in == 8'h56)? 32'h664fd145
	         : (byte_in == 8'h57)? 32'hd7bb41f9
	         : (byte_in == 8'h58)? 32'h4443b158
	         : (byte_in == 8'h59)? 32'hf5b721e4
	         : (byte_in == 8'h5a)? 32'h84e07185
	         : (byte_in == 8'h5b)? 32'h3514e139
	         : (byte_in == 8'h5c)? 32'h27aa9020
	         : (byte_in == 8'h5d)? 32'h965e009c
	         : (byte_in == 8'h5e)? 32'he70950fd
	         : (byte_in == 8'h5f)? 32'h56fdc041
	         : (byte_in == 8'h60)? 32'he6660ae5
	         : (byte_in == 8'h61)? 32'h57929a59
	         : (byte_in == 8'h62)? 32'h26c5ca38
	         : (byte_in == 8'h63)? 32'h97315a84
	         : (byte_in == 8'h64)? 32'h858f2b9d
	         : (byte_in == 8'h65)? 32'h347bbb21
	         : (byte_in == 8'h66)? 32'h452ceb40
	         : (byte_in == 8'h67)? 32'hf4d87bfc
	         : (byte_in == 8'h68)? 32'h67208b5d
	         : (byte_in == 8'h69)? 32'hd6d41be1
	         : (byte_in == 8'h6a)? 32'ha7834b80
	         : (byte_in == 8'h6b)? 32'h1677db3c
	         : (byte_in == 8'h6c)? 32'h04c9aa25
	         : (byte_in == 8'h6d)? 32'hb53d3a99
	         : (byte_in == 8'h6e)? 32'hc46a6af8
	         : (byte_in == 8'h6f)? 32'h759efa44
	         : (byte_in == 8'h70)? 32'h94118e2e
	         : (byte_in == 8'h71)? 32'h25e51e92
	         : (byte_in == 8'h72)? 32'h54b24ef3
	         : (byte_in == 8'h73)? 32'he546de4f
	         : (byte_in == 8'h74)? 32'hf7f8af56
	         : (byte_in == 8'h75)? 32'h460c3fea
	         : (byte_in == 8'h76)? 32'h375b6f8b
	         : (byte_in == 8'h77)? 32'h86afff37
	         : (byte_in == 8'h78)? 32'h15570f96
	         : (byte_in == 8'h79)? 32'ha4a39f2a
	         : (byte_in == 8'h7a)? 32'hd5f4cf4b
	         : (byte_in == 8'h7b)? 32'h64005ff7
	         : (byte_in == 8'h7c)? 32'h76be2eee
	         : (byte_in == 8'h7d)? 32'hc74abe52
	         : (byte_in == 8'h7e)? 32'hb61dee33
	         : (byte_in == 8'h7f)? 32'h07e97e8f
	         : (byte_in == 8'h80)? 32'h44100618
	         : (byte_in == 8'h81)? 32'hf5e496a4
	         : (byte_in == 8'h82)? 32'h84b3c6c5
	         : (byte_in == 8'h83)? 32'h35475679
	         : (byte_in == 8'h84)? 32'h27f92760
	         : (byte_in == 8'h85)? 32'h960db7dc
	         : (byte_in == 8'h86)? 32'he75ae7bd
	         : (byte_in == 8'h87)? 32'h56ae7701
	         : (byte_in == 8'h88)? 32'hc55687a0
	         : (byte_in == 8'h89)? 32'h74a2171c
	         : (byte_in == 8'h8a)? 32'h05f5477d
	         : (byte_in == 8'h8b)? 32'hb401d7c1
	         : (byte_in == 8'h8c)? 32'ha6bfa6d8
	         : (byte_in == 8'h8d)? 32'h174b3664
	         : (byte_in == 8'h8e)? 32'h661c6605
	         : (byte_in == 8'h8f)? 32'hd7e8f6b9
	         : (byte_in == 8'h90)? 32'h366782d3
	         : (byte_in == 8'h91)? 32'h8793126f
	         : (byte_in == 8'h92)? 32'hf6c4420e
	         : (byte_in == 8'h93)? 32'h4730d2b2
	         : (byte_in == 8'h94)? 32'h558ea3ab
	         : (byte_in == 8'h95)? 32'he47a3317
	         : (byte_in == 8'h96)? 32'h952d6376
	         : (byte_in == 8'h97)? 32'h24d9f3ca
	         : (byte_in == 8'h98)? 32'hb721036b
	         : (byte_in == 8'h99)? 32'h06d593d7
	         : (byte_in == 8'h9a)? 32'h7782c3b6
	         : (byte_in == 8'h9b)? 32'hc676530a
	         : (byte_in == 8'h9c)? 32'hd4c82213
	         : (byte_in == 8'h9d)? 32'h653cb2af
	         : (byte_in == 8'h9e)? 32'h146be2ce
	         : (byte_in == 8'h9f)? 32'ha59f7272
	         : (byte_in == 8'ha0)? 32'h1504b8d6
	         : (byte_in == 8'ha1)? 32'ha4f0286a
	         : (byte_in == 8'ha2)? 32'hd5a7780b
	         : (byte_in == 8'ha3)? 32'h6453e8b7
	         : (byte_in == 8'ha4)? 32'h76ed99ae
	         : (byte_in == 8'ha5)? 32'hc7190912
	         : (byte_in == 8'ha6)? 32'hb64e5973
	         : (byte_in == 8'ha7)? 32'h07bac9cf
	         : (byte_in == 8'ha8)? 32'h9442396e
	         : (byte_in == 8'ha9)? 32'h25b6a9d2
	         : (byte_in == 8'haa)? 32'h54e1f9b3
	         : (byte_in == 8'hab)? 32'he515690f
	         : (byte_in == 8'hac)? 32'hf7ab1816
	         : (byte_in == 8'had)? 32'h465f88aa
	         : (byte_in == 8'hae)? 32'h3708d8cb
	         : (byte_in == 8'haf)? 32'h86fc4877
	         : (byte_in == 8'hb0)? 32'h67733c1d
	         : (byte_in == 8'hb1)? 32'hd687aca1
	         : (byte_in == 8'hb2)? 32'ha7d0fcc0
	         : (byte_in == 8'hb3)? 32'h16246c7c
	         : (byte_in == 8'hb4)? 32'h049a1d65
	         : (byte_in == 8'hb5)? 32'hb56e8dd9
	         : (byte_in == 8'hb6)? 32'hc439ddb8
	         : (byte_in == 8'hb7)? 32'h75cd4d04
	         : (byte_in == 8'hb8)? 32'he635bda5
	         : (byte_in == 8'hb9)? 32'h57c12d19
	         : (byte_in == 8'hba)? 32'h26967d78
	         : (byte_in == 8'hbb)? 32'h9762edc4
	         : (byte_in == 8'hbc)? 32'h85dc9cdd
	         : (byte_in == 8'hbd)? 32'h34280c61
	         : (byte_in == 8'hbe)? 32'h457f5c00
	         : (byte_in == 8'hbf)? 32'hf48bccbc
	         : (byte_in == 8'hc0)? 32'hf362b233
	         : (byte_in == 8'hc1)? 32'h4296228f
	         : (byte_in == 8'hc2)? 32'h33c172ee
	         : (byte_in == 8'hc3)? 32'h8235e252
	         : (byte_in == 8'hc4)? 32'h908b934b
	         : (byte_in == 8'hc5)? 32'h217f03f7
	         : (byte_in == 8'hc6)? 32'h50285396
	         : (byte_in == 8'hc7)? 32'he1dcc32a
	         : (byte_in == 8'hc8)? 32'h7224338b
	         : (byte_in == 8'hc9)? 32'hc3d0a337
	         : (byte_in == 8'hca)? 32'hb287f356
	         : (byte_in == 8'hcb)? 32'h037363ea
	         : (byte_in == 8'hcc)? 32'h11cd12f3
	         : (byte_in == 8'hcd)? 32'ha039824f
	         : (byte_in == 8'hce)? 32'hd16ed22e
	         : (byte_in == 8'hcf)? 32'h609a4292
	         : (byte_in == 8'hd0)? 32'h811536f8
	         : (byte_in == 8'hd1)? 32'h30e1a644
	         : (byte_in == 8'hd2)? 32'h41b6f625
	         : (byte_in == 8'hd3)? 32'hf0426699
	         : (byte_in == 8'hd4)? 32'he2fc1780
	         : (byte_in == 8'hd5)? 32'h5308873c
	         : (byte_in == 8'hd6)? 32'h225fd75d
	         : (byte_in == 8'hd7)? 32'h93ab47e1
	         : (byte_in == 8'hd8)? 32'h0053b740
	         : (byte_in == 8'hd9)? 32'hb1a727fc
	         : (byte_in == 8'hda)? 32'hc0f0779d
	         : (byte_in == 8'hdb)? 32'h7104e721
	         : (byte_in == 8'hdc)? 32'h63ba9638
	         : (byte_in == 8'hdd)? 32'hd24e0684
	         : (byte_in == 8'hde)? 32'ha31956e5
	         : (byte_in == 8'hdf)? 32'h12edc659
	         : (byte_in == 8'he0)? 32'ha2760cfd
	         : (byte_in == 8'he1)? 32'h13829c41
	         : (byte_in == 8'he2)? 32'h62d5cc20
	         : (byte_in == 8'he3)? 32'hd3215c9c
	         : (byte_in == 8'he4)? 32'hc19f2d85
	         : (byte_in == 8'he5)? 32'h706bbd39
	         : (byte_in == 8'he6)? 32'h013ced58
	         : (byte_in == 8'he7)? 32'hb0c87de4
	         : (byte_in == 8'he8)? 32'h23308d45
	         : (byte_in == 8'he9)? 32'h92c41df9
	         : (byte_in == 8'hea)? 32'he3934d98
	         : (byte_in == 8'heb)? 32'h5267dd24
	         : (byte_in == 8'hec)? 32'h40d9ac3d
	         : (byte_in == 8'hed)? 32'hf12d3c81
	         : (byte_in == 8'hee)? 32'h807a6ce0
	         : (byte_in == 8'hef)? 32'h318efc5c
	         : (byte_in == 8'hf0)? 32'hd0018836
	         : (byte_in == 8'hf1)? 32'h61f5188a
	         : (byte_in == 8'hf2)? 32'h10a248eb
	         : (byte_in == 8'hf3)? 32'ha156d857
	         : (byte_in == 8'hf4)? 32'hb3e8a94e
	         : (byte_in == 8'hf5)? 32'h021c39f2
	         : (byte_in == 8'hf6)? 32'h734b6993
	         : (byte_in == 8'hf7)? 32'hc2bff92f
	         : (byte_in == 8'hf8)? 32'h5147098e
	         : (byte_in == 8'hf9)? 32'he0b39932
	         : (byte_in == 8'hfa)? 32'h91e4c953
	         : (byte_in == 8'hfb)? 32'h201059ef
	         : (byte_in == 8'hfc)? 32'h32ae28f6
	         : (byte_in == 8'hfd)? 32'h835ab84a
	         : (byte_in == 8'hfe)? 32'hf20de82b
	         :                     32'h43f97897;

endmodule
//}}}

module TABLE30(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'h6ee56854
	         : (byte_in == 8'h02)? 32'h88210c30
	         : (byte_in == 8'h03)? 32'he6c46464
	         : (byte_in == 8'h04)? 32'h3bf3ab2c
	         : (byte_in == 8'h05)? 32'h5516c378
	         : (byte_in == 8'h06)? 32'hb3d2a71c
	         : (byte_in == 8'h07)? 32'hdd37cf48
	         : (byte_in == 8'h08)? 32'ha5e7de5a
	         : (byte_in == 8'h09)? 32'hcb02b60e
	         : (byte_in == 8'h0a)? 32'h2dc6d26a
	         : (byte_in == 8'h0b)? 32'h4323ba3e
	         : (byte_in == 8'h0c)? 32'h9e147576
	         : (byte_in == 8'h0d)? 32'hf0f11d22
	         : (byte_in == 8'h0e)? 32'h16357946
	         : (byte_in == 8'h0f)? 32'h78d01112
	         : (byte_in == 8'h10)? 32'h247febe6
	         : (byte_in == 8'h11)? 32'h4a9a83b2
	         : (byte_in == 8'h12)? 32'hac5ee7d6
	         : (byte_in == 8'h13)? 32'hc2bb8f82
	         : (byte_in == 8'h14)? 32'h1f8c40ca
	         : (byte_in == 8'h15)? 32'h7169289e
	         : (byte_in == 8'h16)? 32'h97ad4cfa
	         : (byte_in == 8'h17)? 32'hf94824ae
	         : (byte_in == 8'h18)? 32'h819835bc
	         : (byte_in == 8'h19)? 32'hef7d5de8
	         : (byte_in == 8'h1a)? 32'h09b9398c
	         : (byte_in == 8'h1b)? 32'h675c51d8
	         : (byte_in == 8'h1c)? 32'hba6b9e90
	         : (byte_in == 8'h1d)? 32'hd48ef6c4
	         : (byte_in == 8'h1e)? 32'h324a92a0
	         : (byte_in == 8'h1f)? 32'h5caffaf4
	         : (byte_in == 8'h20)? 32'hadf2c730
	         : (byte_in == 8'h21)? 32'hc317af64
	         : (byte_in == 8'h22)? 32'h25d3cb00
	         : (byte_in == 8'h23)? 32'h4b36a354
	         : (byte_in == 8'h24)? 32'h96016c1c
	         : (byte_in == 8'h25)? 32'hf8e40448
	         : (byte_in == 8'h26)? 32'h1e20602c
	         : (byte_in == 8'h27)? 32'h70c50878
	         : (byte_in == 8'h28)? 32'h0815196a
	         : (byte_in == 8'h29)? 32'h66f0713e
	         : (byte_in == 8'h2a)? 32'h8034155a
	         : (byte_in == 8'h2b)? 32'heed17d0e
	         : (byte_in == 8'h2c)? 32'h33e6b246
	         : (byte_in == 8'h2d)? 32'h5d03da12
	         : (byte_in == 8'h2e)? 32'hbbc7be76
	         : (byte_in == 8'h2f)? 32'hd522d622
	         : (byte_in == 8'h30)? 32'h898d2cd6
	         : (byte_in == 8'h31)? 32'he7684482
	         : (byte_in == 8'h32)? 32'h01ac20e6
	         : (byte_in == 8'h33)? 32'h6f4948b2
	         : (byte_in == 8'h34)? 32'hb27e87fa
	         : (byte_in == 8'h35)? 32'hdc9befae
	         : (byte_in == 8'h36)? 32'h3a5f8bca
	         : (byte_in == 8'h37)? 32'h54bae39e
	         : (byte_in == 8'h38)? 32'h2c6af28c
	         : (byte_in == 8'h39)? 32'h428f9ad8
	         : (byte_in == 8'h3a)? 32'ha44bfebc
	         : (byte_in == 8'h3b)? 32'hcaae96e8
	         : (byte_in == 8'h3c)? 32'h179959a0
	         : (byte_in == 8'h3d)? 32'h797c31f4
	         : (byte_in == 8'h3e)? 32'h9fb85590
	         : (byte_in == 8'h3f)? 32'hf15d3dc4
	         : (byte_in == 8'h40)? 32'h1b666a73
	         : (byte_in == 8'h41)? 32'h75830227
	         : (byte_in == 8'h42)? 32'h93476643
	         : (byte_in == 8'h43)? 32'hfda20e17
	         : (byte_in == 8'h44)? 32'h2095c15f
	         : (byte_in == 8'h45)? 32'h4e70a90b
	         : (byte_in == 8'h46)? 32'ha8b4cd6f
	         : (byte_in == 8'h47)? 32'hc651a53b
	         : (byte_in == 8'h48)? 32'hbe81b429
	         : (byte_in == 8'h49)? 32'hd064dc7d
	         : (byte_in == 8'h4a)? 32'h36a0b819
	         : (byte_in == 8'h4b)? 32'h5845d04d
	         : (byte_in == 8'h4c)? 32'h85721f05
	         : (byte_in == 8'h4d)? 32'heb977751
	         : (byte_in == 8'h4e)? 32'h0d531335
	         : (byte_in == 8'h4f)? 32'h63b67b61
	         : (byte_in == 8'h50)? 32'h3f198195
	         : (byte_in == 8'h51)? 32'h51fce9c1
	         : (byte_in == 8'h52)? 32'hb7388da5
	         : (byte_in == 8'h53)? 32'hd9dde5f1
	         : (byte_in == 8'h54)? 32'h04ea2ab9
	         : (byte_in == 8'h55)? 32'h6a0f42ed
	         : (byte_in == 8'h56)? 32'h8ccb2689
	         : (byte_in == 8'h57)? 32'he22e4edd
	         : (byte_in == 8'h58)? 32'h9afe5fcf
	         : (byte_in == 8'h59)? 32'hf41b379b
	         : (byte_in == 8'h5a)? 32'h12df53ff
	         : (byte_in == 8'h5b)? 32'h7c3a3bab
	         : (byte_in == 8'h5c)? 32'ha10df4e3
	         : (byte_in == 8'h5d)? 32'hcfe89cb7
	         : (byte_in == 8'h5e)? 32'h292cf8d3
	         : (byte_in == 8'h5f)? 32'h47c99087
	         : (byte_in == 8'h60)? 32'hb694ad43
	         : (byte_in == 8'h61)? 32'hd871c517
	         : (byte_in == 8'h62)? 32'h3eb5a173
	         : (byte_in == 8'h63)? 32'h5050c927
	         : (byte_in == 8'h64)? 32'h8d67066f
	         : (byte_in == 8'h65)? 32'he3826e3b
	         : (byte_in == 8'h66)? 32'h05460a5f
	         : (byte_in == 8'h67)? 32'h6ba3620b
	         : (byte_in == 8'h68)? 32'h13737319
	         : (byte_in == 8'h69)? 32'h7d961b4d
	         : (byte_in == 8'h6a)? 32'h9b527f29
	         : (byte_in == 8'h6b)? 32'hf5b7177d
	         : (byte_in == 8'h6c)? 32'h2880d835
	         : (byte_in == 8'h6d)? 32'h4665b061
	         : (byte_in == 8'h6e)? 32'ha0a1d405
	         : (byte_in == 8'h6f)? 32'hce44bc51
	         : (byte_in == 8'h70)? 32'h92eb46a5
	         : (byte_in == 8'h71)? 32'hfc0e2ef1
	         : (byte_in == 8'h72)? 32'h1aca4a95
	         : (byte_in == 8'h73)? 32'h742f22c1
	         : (byte_in == 8'h74)? 32'ha918ed89
	         : (byte_in == 8'h75)? 32'hc7fd85dd
	         : (byte_in == 8'h76)? 32'h2139e1b9
	         : (byte_in == 8'h77)? 32'h4fdc89ed
	         : (byte_in == 8'h78)? 32'h370c98ff
	         : (byte_in == 8'h79)? 32'h59e9f0ab
	         : (byte_in == 8'h7a)? 32'hbf2d94cf
	         : (byte_in == 8'h7b)? 32'hd1c8fc9b
	         : (byte_in == 8'h7c)? 32'h0cff33d3
	         : (byte_in == 8'h7d)? 32'h621a5b87
	         : (byte_in == 8'h7e)? 32'h84de3fe3
	         : (byte_in == 8'h7f)? 32'hea3b57b7
	         : (byte_in == 8'h80)? 32'hbdd9f5e5
	         : (byte_in == 8'h81)? 32'hd33c9db1
	         : (byte_in == 8'h82)? 32'h35f8f9d5
	         : (byte_in == 8'h83)? 32'h5b1d9181
	         : (byte_in == 8'h84)? 32'h862a5ec9
	         : (byte_in == 8'h85)? 32'he8cf369d
	         : (byte_in == 8'h86)? 32'h0e0b52f9
	         : (byte_in == 8'h87)? 32'h60ee3aad
	         : (byte_in == 8'h88)? 32'h183e2bbf
	         : (byte_in == 8'h89)? 32'h76db43eb
	         : (byte_in == 8'h8a)? 32'h901f278f
	         : (byte_in == 8'h8b)? 32'hfefa4fdb
	         : (byte_in == 8'h8c)? 32'h23cd8093
	         : (byte_in == 8'h8d)? 32'h4d28e8c7
	         : (byte_in == 8'h8e)? 32'habec8ca3
	         : (byte_in == 8'h8f)? 32'hc509e4f7
	         : (byte_in == 8'h90)? 32'h99a61e03
	         : (byte_in == 8'h91)? 32'hf7437657
	         : (byte_in == 8'h92)? 32'h11871233
	         : (byte_in == 8'h93)? 32'h7f627a67
	         : (byte_in == 8'h94)? 32'ha255b52f
	         : (byte_in == 8'h95)? 32'hccb0dd7b
	         : (byte_in == 8'h96)? 32'h2a74b91f
	         : (byte_in == 8'h97)? 32'h4491d14b
	         : (byte_in == 8'h98)? 32'h3c41c059
	         : (byte_in == 8'h99)? 32'h52a4a80d
	         : (byte_in == 8'h9a)? 32'hb460cc69
	         : (byte_in == 8'h9b)? 32'hda85a43d
	         : (byte_in == 8'h9c)? 32'h07b26b75
	         : (byte_in == 8'h9d)? 32'h69570321
	         : (byte_in == 8'h9e)? 32'h8f936745
	         : (byte_in == 8'h9f)? 32'he1760f11
	         : (byte_in == 8'ha0)? 32'h102b32d5
	         : (byte_in == 8'ha1)? 32'h7ece5a81
	         : (byte_in == 8'ha2)? 32'h980a3ee5
	         : (byte_in == 8'ha3)? 32'hf6ef56b1
	         : (byte_in == 8'ha4)? 32'h2bd899f9
	         : (byte_in == 8'ha5)? 32'h453df1ad
	         : (byte_in == 8'ha6)? 32'ha3f995c9
	         : (byte_in == 8'ha7)? 32'hcd1cfd9d
	         : (byte_in == 8'ha8)? 32'hb5ccec8f
	         : (byte_in == 8'ha9)? 32'hdb2984db
	         : (byte_in == 8'haa)? 32'h3dede0bf
	         : (byte_in == 8'hab)? 32'h530888eb
	         : (byte_in == 8'hac)? 32'h8e3f47a3
	         : (byte_in == 8'had)? 32'he0da2ff7
	         : (byte_in == 8'hae)? 32'h061e4b93
	         : (byte_in == 8'haf)? 32'h68fb23c7
	         : (byte_in == 8'hb0)? 32'h3454d933
	         : (byte_in == 8'hb1)? 32'h5ab1b167
	         : (byte_in == 8'hb2)? 32'hbc75d503
	         : (byte_in == 8'hb3)? 32'hd290bd57
	         : (byte_in == 8'hb4)? 32'h0fa7721f
	         : (byte_in == 8'hb5)? 32'h61421a4b
	         : (byte_in == 8'hb6)? 32'h87867e2f
	         : (byte_in == 8'hb7)? 32'he963167b
	         : (byte_in == 8'hb8)? 32'h91b30769
	         : (byte_in == 8'hb9)? 32'hff566f3d
	         : (byte_in == 8'hba)? 32'h19920b59
	         : (byte_in == 8'hbb)? 32'h7777630d
	         : (byte_in == 8'hbc)? 32'haa40ac45
	         : (byte_in == 8'hbd)? 32'hc4a5c411
	         : (byte_in == 8'hbe)? 32'h2261a075
	         : (byte_in == 8'hbf)? 32'h4c84c821
	         : (byte_in == 8'hc0)? 32'ha6bf9f96
	         : (byte_in == 8'hc1)? 32'hc85af7c2
	         : (byte_in == 8'hc2)? 32'h2e9e93a6
	         : (byte_in == 8'hc3)? 32'h407bfbf2
	         : (byte_in == 8'hc4)? 32'h9d4c34ba
	         : (byte_in == 8'hc5)? 32'hf3a95cee
	         : (byte_in == 8'hc6)? 32'h156d388a
	         : (byte_in == 8'hc7)? 32'h7b8850de
	         : (byte_in == 8'hc8)? 32'h035841cc
	         : (byte_in == 8'hc9)? 32'h6dbd2998
	         : (byte_in == 8'hca)? 32'h8b794dfc
	         : (byte_in == 8'hcb)? 32'he59c25a8
	         : (byte_in == 8'hcc)? 32'h38abeae0
	         : (byte_in == 8'hcd)? 32'h564e82b4
	         : (byte_in == 8'hce)? 32'hb08ae6d0
	         : (byte_in == 8'hcf)? 32'hde6f8e84
	         : (byte_in == 8'hd0)? 32'h82c07470
	         : (byte_in == 8'hd1)? 32'hec251c24
	         : (byte_in == 8'hd2)? 32'h0ae17840
	         : (byte_in == 8'hd3)? 32'h64041014
	         : (byte_in == 8'hd4)? 32'hb933df5c
	         : (byte_in == 8'hd5)? 32'hd7d6b708
	         : (byte_in == 8'hd6)? 32'h3112d36c
	         : (byte_in == 8'hd7)? 32'h5ff7bb38
	         : (byte_in == 8'hd8)? 32'h2727aa2a
	         : (byte_in == 8'hd9)? 32'h49c2c27e
	         : (byte_in == 8'hda)? 32'haf06a61a
	         : (byte_in == 8'hdb)? 32'hc1e3ce4e
	         : (byte_in == 8'hdc)? 32'h1cd40106
	         : (byte_in == 8'hdd)? 32'h72316952
	         : (byte_in == 8'hde)? 32'h94f50d36
	         : (byte_in == 8'hdf)? 32'hfa106562
	         : (byte_in == 8'he0)? 32'h0b4d58a6
	         : (byte_in == 8'he1)? 32'h65a830f2
	         : (byte_in == 8'he2)? 32'h836c5496
	         : (byte_in == 8'he3)? 32'hed893cc2
	         : (byte_in == 8'he4)? 32'h30bef38a
	         : (byte_in == 8'he5)? 32'h5e5b9bde
	         : (byte_in == 8'he6)? 32'hb89fffba
	         : (byte_in == 8'he7)? 32'hd67a97ee
	         : (byte_in == 8'he8)? 32'haeaa86fc
	         : (byte_in == 8'he9)? 32'hc04feea8
	         : (byte_in == 8'hea)? 32'h268b8acc
	         : (byte_in == 8'heb)? 32'h486ee298
	         : (byte_in == 8'hec)? 32'h95592dd0
	         : (byte_in == 8'hed)? 32'hfbbc4584
	         : (byte_in == 8'hee)? 32'h1d7821e0
	         : (byte_in == 8'hef)? 32'h739d49b4
	         : (byte_in == 8'hf0)? 32'h2f32b340
	         : (byte_in == 8'hf1)? 32'h41d7db14
	         : (byte_in == 8'hf2)? 32'ha713bf70
	         : (byte_in == 8'hf3)? 32'hc9f6d724
	         : (byte_in == 8'hf4)? 32'h14c1186c
	         : (byte_in == 8'hf5)? 32'h7a247038
	         : (byte_in == 8'hf6)? 32'h9ce0145c
	         : (byte_in == 8'hf7)? 32'hf2057c08
	         : (byte_in == 8'hf8)? 32'h8ad56d1a
	         : (byte_in == 8'hf9)? 32'he430054e
	         : (byte_in == 8'hfa)? 32'h02f4612a
	         : (byte_in == 8'hfb)? 32'h6c11097e
	         : (byte_in == 8'hfc)? 32'hb126c636
	         : (byte_in == 8'hfd)? 32'hdfc3ae62
	         : (byte_in == 8'hfe)? 32'h3907ca06
	         :                     32'h57e2a252;

endmodule
//}}}

module TABLE31(
	byte_in,
	table_out
);

//{{{
input  [7:0]  byte_in;
output [31:0] table_out;

assign table_out = (byte_in == 8'h00)? 32'h00000000
	         : (byte_in == 8'h01)? 32'hd0f4af61
	         : (byte_in == 8'h02)? 32'hce122df3
	         : (byte_in == 8'h03)? 32'h1ee68292
	         : (byte_in == 8'h04)? 32'ha1ec5ec1
	         : (byte_in == 8'h05)? 32'h7118f1a0
	         : (byte_in == 8'h06)? 32'h6ffe7332
	         : (byte_in == 8'h07)? 32'hbf0adc53
	         : (byte_in == 8'h08)? 32'h9c255be5
	         : (byte_in == 8'h09)? 32'h4cd1f484
	         : (byte_in == 8'h0a)? 32'h52377616
	         : (byte_in == 8'h0b)? 32'h82c3d977
	         : (byte_in == 8'h0c)? 32'h3dc90524
	         : (byte_in == 8'h0d)? 32'hed3daa45
	         : (byte_in == 8'h0e)? 32'hf3db28d7
	         : (byte_in == 8'h0f)? 32'h232f87b6
	         : (byte_in == 8'h10)? 32'h1041003e
	         : (byte_in == 8'h11)? 32'hc0b5af5f
	         : (byte_in == 8'h12)? 32'hde532dcd
	         : (byte_in == 8'h13)? 32'h0ea782ac
	         : (byte_in == 8'h14)? 32'hb1ad5eff
	         : (byte_in == 8'h15)? 32'h6159f19e
	         : (byte_in == 8'h16)? 32'h7fbf730c
	         : (byte_in == 8'h17)? 32'haf4bdc6d
	         : (byte_in == 8'h18)? 32'h8c645bdb
	         : (byte_in == 8'h19)? 32'h5c90f4ba
	         : (byte_in == 8'h1a)? 32'h42767628
	         : (byte_in == 8'h1b)? 32'h9282d949
	         : (byte_in == 8'h1c)? 32'h2d88051a
	         : (byte_in == 8'h1d)? 32'hfd7caa7b
	         : (byte_in == 8'h1e)? 32'he39a28e9
	         : (byte_in == 8'h1f)? 32'h336e8788
	         : (byte_in == 8'h20)? 32'hde77cc4c
	         : (byte_in == 8'h21)? 32'h0e83632d
	         : (byte_in == 8'h22)? 32'h1065e1bf
	         : (byte_in == 8'h23)? 32'hc0914ede
	         : (byte_in == 8'h24)? 32'h7f9b928d
	         : (byte_in == 8'h25)? 32'haf6f3dec
	         : (byte_in == 8'h26)? 32'hb189bf7e
	         : (byte_in == 8'h27)? 32'h617d101f
	         : (byte_in == 8'h28)? 32'h425297a9
	         : (byte_in == 8'h29)? 32'h92a638c8
	         : (byte_in == 8'h2a)? 32'h8c40ba5a
	         : (byte_in == 8'h2b)? 32'h5cb4153b
	         : (byte_in == 8'h2c)? 32'he3bec968
	         : (byte_in == 8'h2d)? 32'h334a6609
	         : (byte_in == 8'h2e)? 32'h2dace49b
	         : (byte_in == 8'h2f)? 32'hfd584bfa
	         : (byte_in == 8'h30)? 32'hce36cc72
	         : (byte_in == 8'h31)? 32'h1ec26313
	         : (byte_in == 8'h32)? 32'h0024e181
	         : (byte_in == 8'h33)? 32'hd0d04ee0
	         : (byte_in == 8'h34)? 32'h6fda92b3
	         : (byte_in == 8'h35)? 32'hbf2e3dd2
	         : (byte_in == 8'h36)? 32'ha1c8bf40
	         : (byte_in == 8'h37)? 32'h713c1021
	         : (byte_in == 8'h38)? 32'h52139797
	         : (byte_in == 8'h39)? 32'h82e738f6
	         : (byte_in == 8'h3a)? 32'h9c01ba64
	         : (byte_in == 8'h3b)? 32'h4cf51505
	         : (byte_in == 8'h3c)? 32'hf3ffc956
	         : (byte_in == 8'h3d)? 32'h230b6637
	         : (byte_in == 8'h3e)? 32'h3dede4a5
	         : (byte_in == 8'h3f)? 32'hed194bc4
	         : (byte_in == 8'h40)? 32'h731ebdc2
	         : (byte_in == 8'h41)? 32'ha3ea12a3
	         : (byte_in == 8'h42)? 32'hbd0c9031
	         : (byte_in == 8'h43)? 32'h6df83f50
	         : (byte_in == 8'h44)? 32'hd2f2e303
	         : (byte_in == 8'h45)? 32'h02064c62
	         : (byte_in == 8'h46)? 32'h1ce0cef0
	         : (byte_in == 8'h47)? 32'hcc146191
	         : (byte_in == 8'h48)? 32'hef3be627
	         : (byte_in == 8'h49)? 32'h3fcf4946
	         : (byte_in == 8'h4a)? 32'h2129cbd4
	         : (byte_in == 8'h4b)? 32'hf1dd64b5
	         : (byte_in == 8'h4c)? 32'h4ed7b8e6
	         : (byte_in == 8'h4d)? 32'h9e231787
	         : (byte_in == 8'h4e)? 32'h80c59515
	         : (byte_in == 8'h4f)? 32'h50313a74
	         : (byte_in == 8'h50)? 32'h635fbdfc
	         : (byte_in == 8'h51)? 32'hb3ab129d
	         : (byte_in == 8'h52)? 32'had4d900f
	         : (byte_in == 8'h53)? 32'h7db93f6e
	         : (byte_in == 8'h54)? 32'hc2b3e33d
	         : (byte_in == 8'h55)? 32'h12474c5c
	         : (byte_in == 8'h56)? 32'h0ca1cece
	         : (byte_in == 8'h57)? 32'hdc5561af
	         : (byte_in == 8'h58)? 32'hff7ae619
	         : (byte_in == 8'h59)? 32'h2f8e4978
	         : (byte_in == 8'h5a)? 32'h3168cbea
	         : (byte_in == 8'h5b)? 32'he19c648b
	         : (byte_in == 8'h5c)? 32'h5e96b8d8
	         : (byte_in == 8'h5d)? 32'h8e6217b9
	         : (byte_in == 8'h5e)? 32'h9084952b
	         : (byte_in == 8'h5f)? 32'h40703a4a
	         : (byte_in == 8'h60)? 32'had69718e
	         : (byte_in == 8'h61)? 32'h7d9ddeef
	         : (byte_in == 8'h62)? 32'h637b5c7d
	         : (byte_in == 8'h63)? 32'hb38ff31c
	         : (byte_in == 8'h64)? 32'h0c852f4f
	         : (byte_in == 8'h65)? 32'hdc71802e
	         : (byte_in == 8'h66)? 32'hc29702bc
	         : (byte_in == 8'h67)? 32'h1263addd
	         : (byte_in == 8'h68)? 32'h314c2a6b
	         : (byte_in == 8'h69)? 32'he1b8850a
	         : (byte_in == 8'h6a)? 32'hff5e0798
	         : (byte_in == 8'h6b)? 32'h2faaa8f9
	         : (byte_in == 8'h6c)? 32'h90a074aa
	         : (byte_in == 8'h6d)? 32'h4054dbcb
	         : (byte_in == 8'h6e)? 32'h5eb25959
	         : (byte_in == 8'h6f)? 32'h8e46f638
	         : (byte_in == 8'h70)? 32'hbd2871b0
	         : (byte_in == 8'h71)? 32'h6ddcded1
	         : (byte_in == 8'h72)? 32'h733a5c43
	         : (byte_in == 8'h73)? 32'ha3cef322
	         : (byte_in == 8'h74)? 32'h1cc42f71
	         : (byte_in == 8'h75)? 32'hcc308010
	         : (byte_in == 8'h76)? 32'hd2d60282
	         : (byte_in == 8'h77)? 32'h0222ade3
	         : (byte_in == 8'h78)? 32'h210d2a55
	         : (byte_in == 8'h79)? 32'hf1f98534
	         : (byte_in == 8'h7a)? 32'hef1f07a6
	         : (byte_in == 8'h7b)? 32'h3feba8c7
	         : (byte_in == 8'h7c)? 32'h80e17494
	         : (byte_in == 8'h7d)? 32'h5015dbf5
	         : (byte_in == 8'h7e)? 32'h4ef35967
	         : (byte_in == 8'h7f)? 32'h9e07f606
	         : (byte_in == 8'h80)? 32'h5ad2e31d
	         : (byte_in == 8'h81)? 32'h8a264c7c
	         : (byte_in == 8'h82)? 32'h94c0ceee
	         : (byte_in == 8'h83)? 32'h4434618f
	         : (byte_in == 8'h84)? 32'hfb3ebddc
	         : (byte_in == 8'h85)? 32'h2bca12bd
	         : (byte_in == 8'h86)? 32'h352c902f
	         : (byte_in == 8'h87)? 32'he5d83f4e
	         : (byte_in == 8'h88)? 32'hc6f7b8f8
	         : (byte_in == 8'h89)? 32'h16031799
	         : (byte_in == 8'h8a)? 32'h08e5950b
	         : (byte_in == 8'h8b)? 32'hd8113a6a
	         : (byte_in == 8'h8c)? 32'h671be639
	         : (byte_in == 8'h8d)? 32'hb7ef4958
	         : (byte_in == 8'h8e)? 32'ha909cbca
	         : (byte_in == 8'h8f)? 32'h79fd64ab
	         : (byte_in == 8'h90)? 32'h4a93e323
	         : (byte_in == 8'h91)? 32'h9a674c42
	         : (byte_in == 8'h92)? 32'h8481ced0
	         : (byte_in == 8'h93)? 32'h547561b1
	         : (byte_in == 8'h94)? 32'heb7fbde2
	         : (byte_in == 8'h95)? 32'h3b8b1283
	         : (byte_in == 8'h96)? 32'h256d9011
	         : (byte_in == 8'h97)? 32'hf5993f70
	         : (byte_in == 8'h98)? 32'hd6b6b8c6
	         : (byte_in == 8'h99)? 32'h064217a7
	         : (byte_in == 8'h9a)? 32'h18a49535
	         : (byte_in == 8'h9b)? 32'hc8503a54
	         : (byte_in == 8'h9c)? 32'h775ae607
	         : (byte_in == 8'h9d)? 32'ha7ae4966
	         : (byte_in == 8'h9e)? 32'hb948cbf4
	         : (byte_in == 8'h9f)? 32'h69bc6495
	         : (byte_in == 8'ha0)? 32'h84a52f51
	         : (byte_in == 8'ha1)? 32'h54518030
	         : (byte_in == 8'ha2)? 32'h4ab702a2
	         : (byte_in == 8'ha3)? 32'h9a43adc3
	         : (byte_in == 8'ha4)? 32'h25497190
	         : (byte_in == 8'ha5)? 32'hf5bddef1
	         : (byte_in == 8'ha6)? 32'heb5b5c63
	         : (byte_in == 8'ha7)? 32'h3baff302
	         : (byte_in == 8'ha8)? 32'h188074b4
	         : (byte_in == 8'ha9)? 32'hc874dbd5
	         : (byte_in == 8'haa)? 32'hd6925947
	         : (byte_in == 8'hab)? 32'h0666f626
	         : (byte_in == 8'hac)? 32'hb96c2a75
	         : (byte_in == 8'had)? 32'h69988514
	         : (byte_in == 8'hae)? 32'h777e0786
	         : (byte_in == 8'haf)? 32'ha78aa8e7
	         : (byte_in == 8'hb0)? 32'h94e42f6f
	         : (byte_in == 8'hb1)? 32'h4410800e
	         : (byte_in == 8'hb2)? 32'h5af6029c
	         : (byte_in == 8'hb3)? 32'h8a02adfd
	         : (byte_in == 8'hb4)? 32'h350871ae
	         : (byte_in == 8'hb5)? 32'he5fcdecf
	         : (byte_in == 8'hb6)? 32'hfb1a5c5d
	         : (byte_in == 8'hb7)? 32'h2beef33c
	         : (byte_in == 8'hb8)? 32'h08c1748a
	         : (byte_in == 8'hb9)? 32'hd835dbeb
	         : (byte_in == 8'hba)? 32'hc6d35979
	         : (byte_in == 8'hbb)? 32'h1627f618
	         : (byte_in == 8'hbc)? 32'ha92d2a4b
	         : (byte_in == 8'hbd)? 32'h79d9852a
	         : (byte_in == 8'hbe)? 32'h673f07b8
	         : (byte_in == 8'hbf)? 32'hb7cba8d9
	         : (byte_in == 8'hc0)? 32'h29cc5edf
	         : (byte_in == 8'hc1)? 32'hf938f1be
	         : (byte_in == 8'hc2)? 32'he7de732c
	         : (byte_in == 8'hc3)? 32'h372adc4d
	         : (byte_in == 8'hc4)? 32'h8820001e
	         : (byte_in == 8'hc5)? 32'h58d4af7f
	         : (byte_in == 8'hc6)? 32'h46322ded
	         : (byte_in == 8'hc7)? 32'h96c6828c
	         : (byte_in == 8'hc8)? 32'hb5e9053a
	         : (byte_in == 8'hc9)? 32'h651daa5b
	         : (byte_in == 8'hca)? 32'h7bfb28c9
	         : (byte_in == 8'hcb)? 32'hab0f87a8
	         : (byte_in == 8'hcc)? 32'h14055bfb
	         : (byte_in == 8'hcd)? 32'hc4f1f49a
	         : (byte_in == 8'hce)? 32'hda177608
	         : (byte_in == 8'hcf)? 32'h0ae3d969
	         : (byte_in == 8'hd0)? 32'h398d5ee1
	         : (byte_in == 8'hd1)? 32'he979f180
	         : (byte_in == 8'hd2)? 32'hf79f7312
	         : (byte_in == 8'hd3)? 32'h276bdc73
	         : (byte_in == 8'hd4)? 32'h98610020
	         : (byte_in == 8'hd5)? 32'h4895af41
	         : (byte_in == 8'hd6)? 32'h56732dd3
	         : (byte_in == 8'hd7)? 32'h868782b2
	         : (byte_in == 8'hd8)? 32'ha5a80504
	         : (byte_in == 8'hd9)? 32'h755caa65
	         : (byte_in == 8'hda)? 32'h6bba28f7
	         : (byte_in == 8'hdb)? 32'hbb4e8796
	         : (byte_in == 8'hdc)? 32'h04445bc5
	         : (byte_in == 8'hdd)? 32'hd4b0f4a4
	         : (byte_in == 8'hde)? 32'hca567636
	         : (byte_in == 8'hdf)? 32'h1aa2d957
	         : (byte_in == 8'he0)? 32'hf7bb9293
	         : (byte_in == 8'he1)? 32'h274f3df2
	         : (byte_in == 8'he2)? 32'h39a9bf60
	         : (byte_in == 8'he3)? 32'he95d1001
	         : (byte_in == 8'he4)? 32'h5657cc52
	         : (byte_in == 8'he5)? 32'h86a36333
	         : (byte_in == 8'he6)? 32'h9845e1a1
	         : (byte_in == 8'he7)? 32'h48b14ec0
	         : (byte_in == 8'he8)? 32'h6b9ec976
	         : (byte_in == 8'he9)? 32'hbb6a6617
	         : (byte_in == 8'hea)? 32'ha58ce485
	         : (byte_in == 8'heb)? 32'h75784be4
	         : (byte_in == 8'hec)? 32'hca7297b7
	         : (byte_in == 8'hed)? 32'h1a8638d6
	         : (byte_in == 8'hee)? 32'h0460ba44
	         : (byte_in == 8'hef)? 32'hd4941525
	         : (byte_in == 8'hf0)? 32'he7fa92ad
	         : (byte_in == 8'hf1)? 32'h370e3dcc
	         : (byte_in == 8'hf2)? 32'h29e8bf5e
	         : (byte_in == 8'hf3)? 32'hf91c103f
	         : (byte_in == 8'hf4)? 32'h4616cc6c
	         : (byte_in == 8'hf5)? 32'h96e2630d
	         : (byte_in == 8'hf6)? 32'h8804e19f
	         : (byte_in == 8'hf7)? 32'h58f04efe
	         : (byte_in == 8'hf8)? 32'h7bdfc948
	         : (byte_in == 8'hf9)? 32'hab2b6629
	         : (byte_in == 8'hfa)? 32'hb5cde4bb
	         : (byte_in == 8'hfb)? 32'h65394bda
	         : (byte_in == 8'hfc)? 32'hda339789
	         : (byte_in == 8'hfd)? 32'h0ac738e8
	         : (byte_in == 8'hfe)? 32'h1421ba7a
	         :                     32'hc4d5151b;

endmodule
//}}}

// vim:fdm=marker
